* NGSPICE file created from Top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

.subckt Top CLK_EXT CLK_PLL CLK_SR Data_SR NMOS1_PS1 NMOS1_PS2 NMOS2_PS1 NMOS2_PS2
+ NMOS_PS3 PMOS1_PS1 PMOS1_PS2 PMOS2_PS1 PMOS2_PS2 PMOS_PS3 RST SIGNAL_OUTPUT VGND
+ VPWR d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5]
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1270_ _0612_ net40 VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__and2_1
X_0985_ Shift_Register_Inst.data_out\[16\] net8 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__and2_1
X_1468_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0191_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.go sky130_fd_sc_hd__dfxtp_1
X_1399_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0011_ _0098_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0770_ Signal_Generator_1_0phase_inst.count\[2\] _0280_ VGND VGND VPWR VPWR _0283_
+ sky130_fd_sc_hd__xor2_1
X_1253_ _0563_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nor2_1
X_1322_ Dead_Time_Generator_inst_3.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__and2b_1
X_1184_ _0554_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
X_0968_ Signal_Generator_2_270phase_inst.count\[2\] _0425_ VGND VGND VPWR VPWR _0432_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0899_ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[2\]
+ Signal_Generator_2_90phase_inst.count\[1\] Signal_Generator_2_90phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or4_2
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0822_ net59 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0684_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[1\]
+ Shift_Register_Inst.shift_state\[0\] VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__and3b_1
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0753_ _0270_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_1305_ _0650_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
X_1236_ net33 net6 VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__or2b_1
X_1098_ _0248_ _0250_ Signal_Generator_2_270phase_inst.count\[5\] VGND VGND VPWR VPWR
+ _0508_ sky130_fd_sc_hd__and3_1
X_1167_ _0553_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1021_ net23 _0459_ _0467_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a211oi_1
X_0805_ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0736_ _0258_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
X_1219_ _0556_ _0562_ _0565_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold41 Signal_Generator_1_180phase_inst.direction VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
Xhold30 _0177_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 Signal_Generator_1_270phase_inst.direction VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1004_ _0454_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
X_0719_ _0215_ _0245_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR PMOS1_PS1 sky130_fd_sc_hd__buf_2
XFILLER_0_41_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ _0443_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1398_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0010_ _0097_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
X_1467_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0190_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1321_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_3.count_dt\[1\]
+ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or2b_1
X_1252_ _0565_ _0571_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__nor2_1
X_1183_ _0554_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
X_0967_ Signal_Generator_2_270phase_inst.count\[2\] _0428_ VGND VGND VPWR VPWR _0431_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0898_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.direction
+ _0363_ _0379_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0821_ _0319_ _0322_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__nor2_1
X_0752_ net1 Shift_Register_Inst.data_out\[16\] _0269_ VGND VGND VPWR VPWR _0270_
+ sky130_fd_sc_hd__mux2_1
X_0683_ _0219_ _0220_ Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ net61 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__a41o_1
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1304_ _0625_ _0626_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__and3_1
X_1235_ _0579_ _0586_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1166_ _0553_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
X_1097_ _0248_ _0506_ Signal_Generator_2_90phase_inst.count\[5\] VGND VGND VPWR VPWR
+ _0507_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1020_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] net16
+ _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__a31o_1
X_0804_ _0299_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0735_ Shift_Register_Inst.data_out\[11\] net1 _0257_ VGND VGND VPWR VPWR _0258_
+ sky130_fd_sc_hd__mux2_1
X_1218_ Signal_Generator_1_0phase_inst.count\[4\] _0558_ _0566_ _0570_ VGND VGND VPWR
+ VPWR _0571_ sky130_fd_sc_hd__o22a_1
X_1149_ _0551_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold42 Shift_Register_Inst.shift_state\[0\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 Dead_Time_Generator_inst_3.count_dt\[4\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 Dead_Time_Generator_inst_1.dt\[3\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _0027_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1003_ _0445_ Shift_Register_Inst.data_out\[17\] NMOS2_PS1_prev VGND VGND VPWR VPWR
+ _0454_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0718_ _0233_ _0219_ Shift_Register_Inst.shift_state\[2\] VGND VGND VPWR VPWR _0246_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput21 net21 VGND VGND VPWR VPWR PMOS1_PS2 sky130_fd_sc_hd__clkbuf_4
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0983_ CLK_PLL CLK_EXT Shift_Register_Inst.data_out\[14\] VGND VGND VPWR VPWR _0443_
+ sky130_fd_sc_hd__mux2_2
XFILLER_0_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1397_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0009_ _0096_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
X_1466_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk net72 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
X_1320_ net74 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__inv_2
X_1182_ _0554_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
X_1251_ _0588_ _0601_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0966_ _0056_ _0429_ _0430_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0897_ Signal_Generator_2_0phase_inst.count\[4\] Signal_Generator_2_0phase_inst.direction
+ _0359_ Signal_Generator_2_0phase_inst.count\[5\] VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o31a_1
X_1449_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0054_ _0148_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0820_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0751_ Shift_Register_Inst.shift_state\[0\] _0216_ Shift_Register_Inst.shift_state\[4\]
+ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__or3b_1
X_0682_ Shift_Register_Inst.shift_state\[2\] VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__buf_2
X_1303_ Dead_Time_Generator_inst_2.count_dt\[1\] _0644_ VGND VGND VPWR VPWR _0649_
+ sky130_fd_sc_hd__xor2_1
X_1096_ Shift_Register_Inst.data_out\[8\] VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__inv_2
X_1234_ _0262_ _0578_ _0573_ _0577_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__o211a_1
X_1165_ _0553_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0949_ _0415_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or3b_1
XFILLER_0_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0803_ _0295_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0734_ _0220_ _0221_ _0219_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__and3b_1
XFILLER_0_1_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1079_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_4.count_dt\[1\]
+ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__or2b_1
X_1217_ _0567_ Signal_Generator_1_90phase_inst.count\[4\] _0568_ _0569_ VGND VGND
+ VPWR VPWR _0570_ sky130_fd_sc_hd__a211o_1
X_1148_ _0551_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold32 Signal_Generator_2_180phase_inst.count\[0\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 _0494_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 Dead_Time_Generator_inst_3.go VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 Signal_Generator_1_270phase_inst.direction VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 Shift_Register_Inst.data_out\[15\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1002_ _0453_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_44_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0717_ Shift_Register_Inst.data_out\[6\] VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__buf_2
XFILLER_0_35_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput22 net22 VGND VGND VPWR VPWR PMOS2_PS1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0982_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0426_ _0442_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1465_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0188_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
X_1396_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0008_ _0095_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1181_ _0554_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
X_1250_ _0589_ _0594_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o21a_1
X_0965_ _0424_ _0429_ Signal_Generator_2_270phase_inst.direction VGND VGND VPWR VPWR
+ _0430_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0896_ net69 _0376_ _0377_ _0361_ _0378_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1448_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0053_ _0147_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1379_ clknet_1_1__leaf_CLK_SR _0158_ _0079_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0750_ _0268_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
X_0681_ Shift_Register_Inst.shift_state\[3\] VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__buf_2
X_1302_ _0648_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_1233_ _0583_ _0584_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1164_ _0481_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__buf_4
X_1095_ net14 VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__inv_2
X_0948_ _0403_ _0414_ _0417_ net62 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0879_ Signal_Generator_2_0phase_inst.count\[1\] Signal_Generator_2_0phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0802_ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[2\] Signal_Generator_1_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0733_ _0256_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
X_1216_ _0242_ _0245_ Signal_Generator_1_180phase_inst.count\[4\] VGND VGND VPWR VPWR
+ _0569_ sky130_fd_sc_hd__and3b_1
XFILLER_0_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1078_ Dead_Time_Generator_inst_4.count_dt\[0\] VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__inv_2
X_1147_ _0551_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold22 _0496_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 Dead_Time_Generator_inst_1.go VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 Signal_Generator_2_0phase_inst.direction VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 Signal_Generator_2_0phase_inst.direction VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 Signal_Generator_2_0phase_inst.count\[0\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1001_ PMOS2_PS1_prev _0448_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0716_ _0244_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput23 net23 VGND VGND VPWR VPWR PMOS2_PS2 sky130_fd_sc_hd__clkbuf_4
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0981_ Signal_Generator_2_270phase_inst.count\[4\] Signal_Generator_2_270phase_inst.direction
+ _0422_ Signal_Generator_2_270phase_inst.count\[5\] VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1395_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0014_ _0094_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.direction sky130_fd_sc_hd__dfstp_2
X_1464_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0187_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
X_1180_ _0554_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
X_0964_ _0428_ _0425_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0895_ Signal_Generator_2_0phase_inst.count\[4\] _0359_ VGND VGND VPWR VPWR _0378_
+ sky130_fd_sc_hd__xnor2_1
X_1447_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0052_ _0146_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1378_ clknet_1_0__leaf_CLK_SR _0157_ _0078_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0680_ _0218_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
X_1301_ _0625_ _0626_ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__and3_1
X_1232_ net33 net3 VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__or2b_1
X_1094_ Signal_Generator_2_0phase_inst.count\[4\] _0498_ _0503_ VGND VGND VPWR VPWR
+ _0504_ sky130_fd_sc_hd__o21ai_1
X_1163_ _0552_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
X_0947_ _0415_ _0416_ _0406_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__a21o_1
X_0878_ net58 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0801_ _0297_ _0304_ _0306_ net63 VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0732_ net1 Shift_Register_Inst.data_out\[10\] _0255_ VGND VGND VPWR VPWR _0256_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1215_ _0241_ Shift_Register_Inst.data_out\[6\] VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nor2_2
X_1146_ _0551_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
X_1077_ Dead_Time_Generator_inst_4.count_dt\[3\] VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__inv_2
Xhold56 Signal_Generator_2_90phase_inst.direction VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 Dead_Time_Generator_inst_1.count_dt\[2\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 Signal_Generator_1_180phase_inst.count\[0\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 Signal_Generator_1_270phase_inst.count\[0\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 net86 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1000_ _0452_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_0_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0715_ _0215_ _0242_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
X_1129_ _0538_ net9 VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR PMOS_PS3 sky130_fd_sc_hd__clkbuf_4
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0980_ Signal_Generator_2_270phase_inst.direction _0439_ _0440_ _0424_ _0441_ VGND
+ VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1394_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0173_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.go sky130_fd_sc_hd__dfxtp_1
X_1463_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk net44 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0963_ Signal_Generator_2_270phase_inst.count\[1\] Signal_Generator_2_270phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0894_ Signal_Generator_2_0phase_inst.count\[4\] _0363_ VGND VGND VPWR VPWR _0377_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_40_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1446_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0051_ _0145_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
X_1377_ clknet_1_0__leaf_CLK_SR _0156_ _0077_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1162_ _0552_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
X_1300_ _0644_ _0646_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__nor2_1
X_1231_ _0008_ _0568_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__nand2_1
X_1093_ Signal_Generator_2_180phase_inst.count\[4\] _0499_ _0500_ _0501_ _0502_ VGND
+ VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0946_ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0877_ _0361_ _0364_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__nor2_1
X_1429_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0041_ _0128_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0731_ Shift_Register_Inst.shift_state\[2\] _0233_ Shift_Register_Inst.shift_state\[3\]
+ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or3b_1
X_0800_ _0300_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1145_ _0551_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
X_1214_ _0245_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__inv_2
X_1076_ net37 Dead_Time_Generator_inst_4.count_dt\[4\] VGND VGND VPWR VPWR _0486_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0929_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0401_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__o31a_2
XFILLER_0_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold24 Signal_Generator_2_270phase_inst.count\[0\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 Signal_Generator_1_180phase_inst.direction VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 Signal_Generator_1_90phase_inst.count\[0\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 Dead_Time_Generator_inst_3.count_dt\[3\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 _0670_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0714_ _0229_ _0219_ Shift_Register_Inst.shift_state\[2\] VGND VGND VPWR VPWR _0243_
+ sky130_fd_sc_hd__or3b_1
X_1128_ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[0\]
+ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[0\]
+ _0248_ _0250_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1059_ _0484_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput25 net25 VGND VGND VPWR VPWR SIGNAL_OUTPUT sky130_fd_sc_hd__buf_6
XFILLER_0_11_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1462_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0185_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.go sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1393_ clknet_1_1__leaf_CLK_SR _0172_ _0093_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_0962_ net49 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
X_0893_ _0373_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or3b_1
X_1445_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0050_ _0144_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1376_ clknet_1_0__leaf_CLK_SR _0155_ _0076_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1092_ Shift_Register_Inst.data_out\[8\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0248_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and3b_1
X_1161_ _0552_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
X_1230_ _0568_ _0580_ _0581_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0945_ _0405_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0876_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__and3_1
X_1428_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0040_ _0127_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_1359_ _0212_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0730_ _0254_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
X_1213_ _0242_ _0245_ Signal_Generator_1_270phase_inst.count\[4\] VGND VGND VPWR VPWR
+ _0566_ sky130_fd_sc_hd__and3_1
X_1075_ _0485_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
X_1144_ _0551_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
X_0928_ Signal_Generator_2_180phase_inst.direction VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__inv_2
X_0859_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o31ai_1
Xhold58 Signal_Generator_2_180phase_inst.direction VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 Shift_Register_Inst.shift_state\[4\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 Dead_Time_Generator_inst_1.count_dt\[4\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 Dead_Time_Generator_inst_1.dt\[3\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
Xhold47 _0189_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0713_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__buf_2
X_1127_ _0531_ _0535_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__a21o_1
X_1058_ _0484_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput15 net15 VGND VGND VPWR VPWR NMOS1_PS1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1392_ clknet_1_1__leaf_CLK_SR _0171_ _0092_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1461_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0184_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0961_ _0424_ _0427_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0892_ _0361_ _0372_ _0375_ net80 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__a22o_1
X_1444_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0056_ _0143_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.direction sky130_fd_sc_hd__dfrtp_4
X_1375_ clknet_1_1__leaf_CLK_SR _0154_ _0075_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1091_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] Signal_Generator_2_270phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__and3_1
X_1160_ _0552_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
X_0944_ _0401_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0875_ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[2\]
+ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and3_1
X_1358_ _0545_ _0549_ _0211_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__and3_1
X_1427_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0039_ _0126_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1289_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_2.count_dt\[1\]
+ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1212_ _0445_ net7 VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2_1
X_1074_ _0485_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1143_ _0551_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
X_0927_ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[2\]
+ Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or4_2
X_0789_ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__and2_1
X_0858_ _0340_ _0347_ _0349_ net68 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold37 Signal_Generator_2_180phase_inst.direction VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
Xhold26 Signal_Generator_2_90phase_inst.count\[0\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 _0621_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 _0005_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 Signal_Generator_1_0phase_inst.count\[4\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0712_ Shift_Register_Inst.data_out\[5\] VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_2
X_1126_ net10 VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__inv_2
X_1057_ _0484_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput16 net16 VGND VGND VPWR VPWR NMOS1_PS2 sky130_fd_sc_hd__buf_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1109_ _0500_ _0516_ _0517_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1391_ clknet_1_1__leaf_CLK_SR _0170_ _0091_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1460_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0183_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0960_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0891_ _0373_ _0374_ _0364_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a21o_1
X_1443_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0048_ _0142_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.count\[5\] sky130_fd_sc_hd__dfstp_1
X_1374_ clknet_1_0__leaf_CLK_SR _0153_ _0074_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ Shift_Register_Inst.data_out\[7\] _0250_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__nor2_1
X_0943_ Signal_Generator_2_180phase_inst.count\[2\] Signal_Generator_2_180phase_inst.count\[1\]
+ Signal_Generator_2_180phase_inst.count\[0\] Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0874_ Signal_Generator_2_0phase_inst.count\[1\] Signal_Generator_2_0phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__and2_1
X_1288_ Dead_Time_Generator_inst_2.count_dt\[0\] VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__inv_2
X_1357_ _0487_ _0207_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__xnor2_1
X_1426_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0038_ _0125_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1142_ _0481_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__buf_4
X_1211_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__inv_2
X_1073_ _0485_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
X_0926_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0384_ _0400_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0857_ _0343_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or2_1
Xhold38 Signal_Generator_1_90phase_inst.direction VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
X_0788_ Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ _0295_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__o31a_1
X_1409_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0021_ _0108_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.direction sky130_fd_sc_hd__dfstp_1
Xhold27 Signal_Generator_1_0phase_inst.count\[0\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold16 Shift_Register_Inst.data_out\[16\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 Dead_Time_Generator_inst_3.count_dt\[2\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0711_ _0240_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_1__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_1125_ _0500_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or4_1
X_1056_ _0484_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
X_0909_ _0382_ _0387_ net65 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a21oi_1
Xoutput17 net17 VGND VGND VPWR VPWR NMOS2_PS1 sky130_fd_sc_hd__clkbuf_4
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1108_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] Signal_Generator_2_180phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1039_ _0262_ net36 _0472_ _0474_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ clknet_1_1__leaf_CLK_SR _0169_ _0090_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0890_ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__a31o_1
X_1442_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0047_ _0141_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.count\[4\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_10_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1373_ clknet_1_1__leaf_CLK_SR _0152_ _0073_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0942_ _0403_ _0410_ _0412_ net62 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__a22o_1
X_0873_ Signal_Generator_2_0phase_inst.count\[5\] Signal_Generator_2_0phase_inst.count\[4\]
+ _0359_ _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o31a_1
X_1425_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0037_ _0124_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_2
X_1287_ Dead_Time_Generator_inst_2.count_dt\[3\] VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__inv_2
X_1356_ _0210_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1141_ _0550_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
X_1210_ _0556_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__nor2_1
X_1072_ _0485_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
X_0925_ Signal_Generator_2_90phase_inst.count\[4\] Signal_Generator_2_90phase_inst.direction
+ _0380_ Signal_Generator_2_90phase_inst.count\[5\] VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__o31a_1
X_0787_ Signal_Generator_1_90phase_inst.direction VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__inv_2
X_0856_ Signal_Generator_1_270phase_inst.count\[2\] _0341_ VGND VGND VPWR VPWR _0348_
+ sky130_fd_sc_hd__xor2_1
Xhold17 _0174_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0034_ _0107_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
Xhold28 Dead_Time_Generator_inst_1.dt\[4\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 Shift_Register_Inst.shift_state\[1\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ _0661_ _0672_ _0660_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0710_ _0215_ Dead_Time_Generator_inst_1.dt\[4\] _0239_ VGND VGND VPWR VPWR _0240_
+ sky130_fd_sc_hd__mux2_1
X_1124_ _0248_ _0250_ Signal_Generator_2_270phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0534_ sky130_fd_sc_hd__and3_1
X_1055_ _0484_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput18 net18 VGND VGND VPWR VPWR NMOS2_PS2 sky130_fd_sc_hd__clkbuf_4
X_0908_ _0386_ _0383_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__or2_1
X_0839_ Signal_Generator_1_180phase_inst.count\[4\] _0317_ VGND VGND VPWR VPWR _0336_
+ sky130_fd_sc_hd__xnor2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1107_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and3_1
X_1038_ _0480_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1441_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0046_ _0140_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.count\[3\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1372_ clknet_1_1__leaf_CLK_SR _0151_ _0072_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0941_ _0406_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0872_ Signal_Generator_2_0phase_inst.direction VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1355_ _0545_ _0549_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__and3_1
X_1424_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0036_ _0123_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1286_ net37 Dead_Time_Generator_inst_2.count_dt\[4\] VGND VGND VPWR VPWR _0633_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1071_ _0485_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1140_ _0497_ _0545_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and3_1
X_0924_ net81 _0397_ _0398_ _0382_ _0399_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a32o_1
X_0786_ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[1\]
+ Signal_Generator_1_90phase_inst.count\[3\] Signal_Generator_1_90phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__or4_2
X_0855_ Signal_Generator_1_270phase_inst.count\[2\] _0344_ VGND VGND VPWR VPWR _0347_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold29 Dead_Time_Generator_inst_1.count_dt\[3\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0033_ _0106_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[4\] sky130_fd_sc_hd__dfstp_2
Xhold18 Dead_Time_Generator_inst_3.count_dt\[0\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ Dead_Time_Generator_inst_3.count_dt\[3\] Dead_Time_Generator_inst_3.count_dt\[2\]
+ Dead_Time_Generator_inst_3.count_dt\[1\] _0669_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__and4_1
X_1269_ Dead_Time_Generator_inst_1.count_dt\[0\] _0612_ net40 VGND VGND VPWR VPWR
+ _0622_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1123_ _0248_ _0250_ Signal_Generator_2_180phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0533_ sky130_fd_sc_hd__and3b_1
X_1054_ _0482_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__buf_4
X_0907_ Signal_Generator_2_90phase_inst.count\[1\] Signal_Generator_2_90phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0838_ Signal_Generator_1_180phase_inst.count\[4\] _0321_ VGND VGND VPWR VPWR _0335_
+ sky130_fd_sc_hd__or2_1
Xoutput19 net19 VGND VGND VPWR VPWR NMOS_PS3 sky130_fd_sc_hd__clkbuf_4
X_0769_ _0014_ _0281_ _0282_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1106_ Shift_Register_Inst.data_out\[8\] Signal_Generator_2_90phase_inst.count\[3\]
+ Shift_Register_Inst.data_out\[7\] VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__and3b_1
XFILLER_0_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1037_ net31 _0477_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1440_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0045_ _0139_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.count\[2\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0001_ _0071_ VGND VGND VPWR
+ VPWR NMOS1_PS2_prev sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ Signal_Generator_2_180phase_inst.count\[2\] _0404_ VGND VGND VPWR VPWR _0411_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0871_ Signal_Generator_2_0phase_inst.count\[3\] Signal_Generator_2_0phase_inst.count\[2\]
+ Signal_Generator_2_0phase_inst.count\[1\] Signal_Generator_2_0phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__or4_2
X_1354_ _0207_ _0208_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__and2b_1
X_1423_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0042_ _0122_ VGND VGND VPWR
+ VPWR Signal_Generator_2_0phase_inst.direction sky130_fd_sc_hd__dfstp_1
X_1285_ _0482_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1070_ _0485_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
X_0923_ Signal_Generator_2_90phase_inst.count\[4\] _0380_ VGND VGND VPWR VPWR _0399_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0854_ _0028_ _0345_ _0346_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a21oi_1
X_0785_ net73 Signal_Generator_1_0phase_inst.direction _0278_ _0294_ VGND VGND VPWR
+ VPWR _0013_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1268_ _0613_ net39 _0618_ _0619_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a221o_1
X_1406_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0032_ _0105_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[3\] sky130_fd_sc_hd__dfstp_1
X_1337_ _0545_ _0549_ _0675_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a21oi_1
Xhold19 _0186_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
X_1199_ _0482_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1122_ _0250_ Signal_Generator_2_90phase_inst.count\[1\] _0248_ VGND VGND VPWR VPWR
+ _0532_ sky130_fd_sc_hd__and3b_1
X_1053_ _0483_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0906_ net51 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__inv_2
X_0837_ _0331_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or3b_1
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0768_ _0276_ _0281_ net75 VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a21oi_1
X_0699_ _0215_ Dead_Time_Generator_inst_1.dt\[1\] _0231_ VGND VGND VPWR VPWR _0232_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1105_ net12 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1036_ _0479_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1019_ net21 _0458_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1370_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0007_ _0070_ VGND VGND VPWR
+ VPWR PMOS2_PS2_prev sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_2__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_0870_ Signal_Generator_1_270phase_inst.count\[4\] net77 _0342_ _0358_ VGND VGND
+ VPWR VPWR _0027_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1422_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk net78 _0121_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[5\] sky130_fd_sc_hd__dfstp_1
X_1284_ _0625_ _0626_ _0631_ net50 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__o2bb2a_1
X_1353_ Dead_Time_Generator_inst_4.count_dt\[1\] _0201_ Dead_Time_Generator_inst_4.count_dt\[2\]
+ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0999_ _0445_ Shift_Register_Inst.data_out\[17\] NMOS1_PS1_prev VGND VGND VPWR VPWR
+ _0452_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ Signal_Generator_2_90phase_inst.count\[4\] _0384_ VGND VGND VPWR VPWR _0398_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0853_ _0340_ _0345_ net68 VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a21oi_1
X_1405_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0031_ _0104_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[2\] sky130_fd_sc_hd__dfstp_2
X_0784_ Signal_Generator_1_0phase_inst.count\[4\] Signal_Generator_1_0phase_inst.direction
+ _0274_ Signal_Generator_1_0phase_inst.count\[5\] VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__o31a_1
X_1198_ _0482_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
X_1267_ Dead_Time_Generator_inst_1.count_dt\[4\] net37 VGND VGND VPWR VPWR _0620_
+ sky130_fd_sc_hd__and2b_1
Xinput1 Data_SR VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_1336_ _0661_ _0672_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1052_ _0483_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
X_1121_ Signal_Generator_2_0phase_inst.count\[1\] _0498_ VGND VGND VPWR VPWR _0531_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0905_ _0382_ _0385_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__nor2_1
X_0836_ _0319_ _0330_ _0333_ net66 VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a22o_1
X_0767_ _0280_ _0277_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0698_ Shift_Register_Inst.shift_state\[4\] _0227_ _0216_ VGND VGND VPWR VPWR _0231_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ net71 VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1035_ net31 _0475_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and2_1
X_1104_ _0511_ _0512_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0819_ Signal_Generator_1_180phase_inst.count\[3\] Signal_Generator_1_180phase_inst.count\[2\]
+ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__and3_1
X_1018_ NMOS2_PS2_prev _0466_ _0456_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0026_ _0120_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_1283_ _0607_ _0611_ _0631_ _0632_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__a211oi_1
X_1352_ Dead_Time_Generator_inst_4.count_dt\[2\] Dead_Time_Generator_inst_4.count_dt\[1\]
+ _0201_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0998_ _0451_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0921_ _0394_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or3b_1
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0783_ Signal_Generator_1_0phase_inst.direction _0291_ _0292_ _0276_ _0293_ VGND
+ VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a32o_1
X_0852_ _0344_ _0341_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1404_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0030_ _0103_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[1\] sky130_fd_sc_hd__dfstp_1
X_1335_ _0545_ _0549_ _0674_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1197_ _0482_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__inv_2
X_1266_ _0614_ Dead_Time_Generator_inst_1.dt\[2\] net39 _0613_ VGND VGND VPWR VPWR
+ _0619_ sky130_fd_sc_hd__o22a_1
Xinput2 RST VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1051_ _0483_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
X_1120_ _0521_ _0527_ _0528_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0904_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0697_ net67 _0228_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__xnor2_1
X_0835_ _0331_ _0332_ _0322_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0766_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1318_ net37 Dead_Time_Generator_inst_3.count_dt\[4\] VGND VGND VPWR VPWR _0659_
+ sky130_fd_sc_hd__or2b_1
X_1249_ _0589_ _0594_ _0595_ _0600_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1034_ _0478_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
X_1103_ net13 _0504_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0818_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0749_ net79 net1 _0267_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1017_ _0445_ Shift_Register_Inst.data_out\[17\] VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1351_ _0206_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
X_1420_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0025_ _0119_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_1282_ _0614_ _0627_ _0613_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0997_ PMOS1_PS2_prev _0448_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0920_ _0382_ _0393_ _0396_ net65 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a22o_1
X_0782_ Signal_Generator_1_0phase_inst.count\[4\] _0274_ VGND VGND VPWR VPWR _0293_
+ sky130_fd_sc_hd__xnor2_1
X_0851_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nor2_1
X_1265_ _0614_ Dead_Time_Generator_inst_1.dt\[2\] _0615_ _0616_ _0617_ VGND VGND VPWR
+ VPWR _0618_ sky130_fd_sc_hd__a221o_1
X_1403_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0029_ _0102_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_1
X_1334_ _0672_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__nand2_1
X_1196_ _0555_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 d1[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_0_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1050_ _0483_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
X_0903_ Signal_Generator_2_90phase_inst.count\[3\] Signal_Generator_2_90phase_inst.count\[2\]
+ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__and3_1
X_0834_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a31o_1
X_0765_ net52 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
X_0696_ _0229_ _0230_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__nand2_1
X_1317_ _0625_ _0626_ _0623_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a21oi_1
X_1248_ _0589_ _0594_ _0595_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o22a_1
X_1179_ _0554_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1102_ _0505_ _0510_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1033_ _0474_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and2_1
X_0817_ Signal_Generator_1_180phase_inst.count\[5\] Signal_Generator_1_180phase_inst.count\[4\]
+ _0317_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o31a_2
XFILLER_0_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0748_ _0219_ _0220_ _0221_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__and3_1
X_0679_ _0215_ Dead_Time_Generator_inst_1.dt\[0\] _0217_ VGND VGND VPWR VPWR _0218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1016_ _0462_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ Dead_Time_Generator_inst_1.count_dt\[3\] Dead_Time_Generator_inst_1.count_dt\[2\]
+ Dead_Time_Generator_inst_1.count_dt\[1\] _0622_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__and4_1
X_1350_ _0545_ _0549_ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__and3_1
X_0996_ _0450_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0850_ net48 VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
X_1402_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0035_ _0101_ VGND VGND VPWR
+ VPWR Signal_Generator_1_90phase_inst.direction sky130_fd_sc_hd__dfstp_1
X_0781_ Signal_Generator_1_0phase_inst.count\[4\] _0278_ VGND VGND VPWR VPWR _0292_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1264_ Dead_Time_Generator_inst_1.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__and2b_1
Xinput4 d1[1] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_1333_ Dead_Time_Generator_inst_3.count_dt\[1\] _0669_ VGND VGND VPWR VPWR _0673_
+ sky130_fd_sc_hd__or2_1
X_1195_ _0555_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__inv_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0979_ Signal_Generator_2_270phase_inst.count\[4\] _0422_ VGND VGND VPWR VPWR _0441_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0902_ Signal_Generator_2_90phase_inst.count\[1\] Signal_Generator_2_90phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__and2_1
X_0833_ _0321_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0764_ _0276_ _0279_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__nor2_1
X_0695_ net61 _0227_ net64 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__o21ai_1
X_1316_ _0658_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
X_1247_ _0568_ _0596_ _0597_ _0598_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__o41a_1
X_1178_ _0554_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
X_1032_ Dead_Time_Generator_inst_4.go net5 _0262_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1101_ _0504_ net13 _0505_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__a2bb2o_1
X_0747_ _0266_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_0816_ Signal_Generator_1_180phase_inst.direction VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0678_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[0\]
+ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__or3_1
Xclkbuf_3_3__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1015_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] net15
+ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _0625_ _0626_ _0630_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ _0445_ Shift_Register_Inst.data_out\[17\] NMOS2_PS2_prev VGND VGND VPWR VPWR
+ _0450_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0780_ _0288_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__or3b_1
X_1401_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0013_ _0100_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_1194_ _0555_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__inv_2
X_1263_ Dead_Time_Generator_inst_1.count_dt\[0\] Dead_Time_Generator_inst_1.dt\[0\]
+ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__and2b_1
Xinput5 d1[2] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_1332_ Dead_Time_Generator_inst_3.count_dt\[1\] _0669_ VGND VGND VPWR VPWR _0672_
+ sky130_fd_sc_hd__nand2_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0978_ Signal_Generator_2_270phase_inst.count\[4\] _0426_ VGND VGND VPWR VPWR _0440_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0901_ Signal_Generator_2_90phase_inst.count\[5\] Signal_Generator_2_90phase_inst.count\[4\]
+ _0380_ _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o31a_1
X_0832_ _0317_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nand2_1
X_0763_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1315_ _0625_ _0626_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0694_ Shift_Register_Inst.shift_state\[1\] _0227_ _0228_ VGND VGND VPWR VPWR _0229_
+ sky130_fd_sc_hd__or3_2
X_1246_ _0242_ _0245_ Signal_Generator_1_0phase_inst.count\[2\] VGND VGND VPWR VPWR
+ _0599_ sky130_fd_sc_hd__or3_1
X_1177_ _0554_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1100_ _0507_ _0508_ _0509_ _0498_ Signal_Generator_2_0phase_inst.count\[5\] VGND
+ VGND VPWR VPWR _0510_ sky130_fd_sc_hd__o32a_1
XFILLER_0_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1031_ _0476_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0746_ net1 net76 _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
X_0815_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[3\] Signal_Generator_1_180phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__or4_2
XFILLER_0_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0677_ Shift_Register_Inst.shift_state\[3\] Shift_Register_Inst.shift_state\[2\]
+ Shift_Register_Inst.shift_state\[1\] VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__or3_2
X_1229_ _0242_ _0245_ Signal_Generator_1_270phase_inst.count\[0\] VGND VGND VPWR VPWR
+ _0582_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1014_ net17 _0456_ _0459_ net22 VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a22o_1
X_0729_ _0215_ Shift_Register_Inst.data_out\[9\] _0253_ VGND VGND VPWR VPWR _0254_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0994_ _0449_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1331_ _0544_ _0548_ _0669_ _0671_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a211oi_1
X_1400_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0012_ _0099_ VGND VGND VPWR
+ VPWR Signal_Generator_1_0phase_inst.count\[4\] sky130_fd_sc_hd__dfrtp_4
X_1193_ _0555_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__inv_2
X_1262_ Dead_Time_Generator_inst_1.dt\[1\] Dead_Time_Generator_inst_1.count_dt\[1\]
+ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or2b_1
Xinput6 d1[3] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0977_ _0436_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or3b_1
XFILLER_0_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ Signal_Generator_2_90phase_inst.direction VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0693_ Shift_Register_Inst.shift_state\[4\] _0216_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__and2_1
X_0831_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ Signal_Generator_1_180phase_inst.count\[2\] Signal_Generator_1_180phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0762_ Signal_Generator_1_0phase_inst.count\[3\] Signal_Generator_1_0phase_inst.count\[2\]
+ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__and3_1
X_1314_ Dead_Time_Generator_inst_2.count_dt\[3\] _0651_ Dead_Time_Generator_inst_2.count_dt\[4\]
+ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a21o_1
Xclkbuf_0_Dead_Time_Generator_inst_1.clk Dead_Time_Generator_inst_1.clk VGND VGND
+ VPWR VPWR clknet_0_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_1245_ _0557_ Signal_Generator_1_90phase_inst.count\[2\] VGND VGND VPWR VPWR _0598_
+ sky130_fd_sc_hd__and2b_1
X_1176_ _0554_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1030_ _0474_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0299_ _0316_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__a31o_1
X_0676_ net1 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0745_ _0259_ _0233_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_1
X_1228_ _0557_ Signal_Generator_1_90phase_inst.count\[0\] _0241_ VGND VGND VPWR VPWR
+ _0581_ sky130_fd_sc_hd__and3b_1
X_1159_ _0552_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1013_ net20 _0458_ Shift_Register_Inst.data_out\[11\] Shift_Register_Inst.data_out\[12\]
+ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a211o_1
X_0728_ _0220_ _0229_ Shift_Register_Inst.shift_state\[3\] VGND VGND VPWR VPWR _0253_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ PMOS2_PS2_prev _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1261_ net70 VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__inv_2
X_1330_ net43 net38 VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nor2_1
X_1192_ _0555_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 d1[4] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_0976_ _0424_ _0435_ _0438_ Signal_Generator_2_270phase_inst.direction VGND VGND
+ VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1459_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0182_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ _0319_ _0326_ _0328_ net66 VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0692_ Shift_Register_Inst.shift_state\[0\] VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__inv_2
X_0761_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__and2_1
X_1313_ _0656_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
X_1244_ _0241_ _0557_ Signal_Generator_1_180phase_inst.count\[2\] VGND VGND VPWR VPWR
+ _0597_ sky130_fd_sc_hd__and3b_1
X_1175_ _0481_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0959_ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[2\]
+ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 d2[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
X_0813_ Signal_Generator_1_90phase_inst.count\[4\] Signal_Generator_1_90phase_inst.direction
+ _0295_ Signal_Generator_1_90phase_inst.count\[5\] VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0744_ _0264_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
X_1158_ _0552_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
X_1227_ _0241_ _0557_ Signal_Generator_1_180phase_inst.count\[0\] VGND VGND VPWR VPWR
+ _0580_ sky130_fd_sc_hd__and3b_1
X_1089_ Shift_Register_Inst.data_out\[7\] Shift_Register_Inst.data_out\[8\] VGND VGND
+ VPWR VPWR _0499_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1012_ net24 _0458_ _0459_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0460_
+ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a221o_2
X_0727_ _0252_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0992_ Shift_Register_Inst.data_out\[16\] Shift_Register_Inst.data_out\[17\] VGND
+ VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or2b_1
XFILLER_0_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput8 d1[5] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
X_1191_ _0555_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1260_ net54 VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ _0436_ _0437_ _0427_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1389_ clknet_1_1__leaf_CLK_SR _0168_ _0089_ VGND VGND VPWR VPWR Shift_Register_Inst.shift_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_1458_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0181_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_4__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ Signal_Generator_1_0phase_inst.count\[5\] Signal_Generator_1_0phase_inst.count\[4\]
+ _0274_ _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__o31a_1
X_0691_ _0226_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
X_1312_ _0625_ _0626_ _0655_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and3_1
X_1243_ _0241_ _0557_ Signal_Generator_1_270phase_inst.count\[2\] VGND VGND VPWR VPWR
+ _0596_ sky130_fd_sc_hd__and3_1
X_1174_ _0553_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
X_0958_ Signal_Generator_2_270phase_inst.count\[1\] Signal_Generator_2_270phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0889_ _0363_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0812_ _0313_ _0314_ _0297_ _0315_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 d2[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_0743_ net1 _0262_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1157_ _0552_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
X_1226_ _0573_ _0577_ net33 _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a211o_1
X_1088_ _0248_ _0250_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1011_ Shift_Register_Inst.data_out\[12\] VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__inv_2
X_0726_ _0215_ _0250_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1209_ Signal_Generator_1_0phase_inst.count\[5\] _0558_ _0560_ _0561_ VGND VGND VPWR
+ VPWR _0562_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0709_ _0238_ _0219_ Shift_Register_Inst.shift_state\[2\] VGND VGND VPWR VPWR _0239_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0991_ _0447_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_0_26_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1474_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0197_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_3.go sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ _0555_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__inv_2
Xinput9 d2[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a31o_1
X_1457_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0180_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_2.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
X_1388_ clknet_1_0__leaf_CLK_SR _0167_ _0088_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0690_ _0222_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1311_ _0634_ _0651_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__xnor2_1
X_1242_ net33 net5 VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or2b_1
X_1173_ _0553_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0957_ Signal_Generator_2_270phase_inst.count\[5\] Signal_Generator_2_270phase_inst.count\[4\]
+ _0422_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o31a_2
X_0888_ _0359_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__nand2_1
X_0811_ Signal_Generator_1_90phase_inst.count\[4\] _0295_ VGND VGND VPWR VPWR _0315_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput12 d2[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_0742_ _0259_ _0229_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__or2_1
X_1156_ _0552_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
X_1225_ net4 VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__inv_2
X_1087_ _0486_ net47 VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] VGND
+ VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and2b_1
X_0725_ _0220_ _0238_ Shift_Register_Inst.shift_state\[3\] VGND VGND VPWR VPWR _0251_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1208_ _0242_ _0312_ _0245_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a21oi_1
X_1139_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0708_ Shift_Register_Inst.shift_state\[1\] Shift_Register_Inst.shift_state\[0\]
+ _0228_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0990_ _0445_ Shift_Register_Inst.data_out\[17\] NMOS1_PS2_prev VGND VGND VPWR VPWR
+ _0447_ sky130_fd_sc_hd__and3_1
X_1473_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0196_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ _0426_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1387_ clknet_1_0__leaf_CLK_SR _0166_ _0087_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_1456_ clknet_1_0__leaf_CLK_SR _0179_ _0150_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ _0654_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_1241_ _0568_ _0590_ _0591_ _0592_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o41a_1
XFILLER_0_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1172_ _0553_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
X_0956_ Signal_Generator_2_270phase_inst.direction VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0887_ Signal_Generator_2_0phase_inst.count\[2\] Signal_Generator_2_0phase_inst.count\[1\]
+ Signal_Generator_2_0phase_inst.count\[0\] Signal_Generator_2_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__o31ai_1
X_1439_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0044_ _0138_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.count\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 d2[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_0_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0810_ Signal_Generator_1_90phase_inst.count\[4\] _0299_ Signal_Generator_1_90phase_inst.direction
+ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0741_ net33 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_4
X_1224_ _0568_ _0574_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__or4_1
X_1155_ _0552_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
X_1086_ _0487_ net39 _0492_ net46 _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__a221o_1
X_0939_ Signal_Generator_2_180phase_inst.count\[2\] _0407_ VGND VGND VPWR VPWR _0410_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0724_ Shift_Register_Inst.data_out\[8\] VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1207_ _0242_ _0245_ Signal_Generator_1_270phase_inst.count\[5\] _0559_ VGND VGND
+ VPWR VPWR _0560_ sky130_fd_sc_hd__a31o_1
X_1069_ _0485_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
X_1138_ _0546_ _0547_ _0530_ _0514_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0707_ _0237_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1472_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0195_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0972_ _0422_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__nand2_1
X_1455_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0178_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[4\] sky130_fd_sc_hd__dfxtp_1
X_1386_ clknet_1_0__leaf_CLK_SR _0165_ _0086_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1240_ _0242_ _0245_ Signal_Generator_1_0phase_inst.count\[3\] VGND VGND VPWR VPWR
+ _0593_ sky130_fd_sc_hd__or3_1
X_1171_ _0553_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0955_ Signal_Generator_2_270phase_inst.count\[3\] Signal_Generator_2_270phase_inst.count\[2\]
+ Signal_Generator_2_270phase_inst.count\[1\] Signal_Generator_2_270phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or4_2
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ _0361_ _0368_ _0370_ net69 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1438_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0043_ _0137_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_1
X_1369_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0003_ _0069_ VGND VGND VPWR
+ VPWR NMOS2_PS2_prev sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput14 d2[5] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_0740_ _0261_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
X_1154_ _0552_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
X_1223_ _0241_ _0557_ Signal_Generator_1_270phase_inst.count\[1\] VGND VGND VPWR VPWR
+ _0576_ sky130_fd_sc_hd__and3_1
X_1085_ Dead_Time_Generator_inst_4.count_dt\[4\] net37 VGND VGND VPWR VPWR _0495_
+ sky130_fd_sc_hd__and2b_1
X_0938_ _0049_ _0408_ _0409_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a21oi_1
X_0869_ Signal_Generator_1_270phase_inst.count\[4\] Signal_Generator_1_270phase_inst.direction
+ _0338_ Signal_Generator_1_270phase_inst.count\[5\] VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0723_ _0249_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1137_ _0540_ _0537_ _0539_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__nand3b_1
X_1206_ _0242_ _0245_ Signal_Generator_1_180phase_inst.count\[5\] VGND VGND VPWR VPWR
+ _0559_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1068_ _0485_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0706_ _0215_ Dead_Time_Generator_inst_1.dt\[3\] _0236_ VGND VGND VPWR VPWR _0237_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1471_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0194_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ Signal_Generator_2_270phase_inst.count\[2\] Signal_Generator_2_270phase_inst.count\[1\]
+ Signal_Generator_2_270phase_inst.count\[0\] Signal_Generator_2_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1454_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk net55 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ clknet_1_0__leaf_CLK_SR _0164_ _0085_ VGND VGND VPWR VPWR Dead_Time_Generator_inst_1.dt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1170_ _0553_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
X_0954_ Signal_Generator_2_180phase_inst.count\[4\] net83 _0405_ _0421_ VGND VGND
+ VPWR VPWR _0048_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0885_ _0364_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__or2_1
X_1437_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0049_ _0136_ VGND VGND VPWR
+ VPWR Signal_Generator_2_180phase_inst.direction sky130_fd_sc_hd__dfstp_1
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1299_ _0635_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__and2_1
X_1368_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk net84 _0068_ VGND VGND VPWR
+ VPWR PMOS1_PS2_prev sky130_fd_sc_hd__dfstp_1
X_1153_ _0481_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__buf_4
X_1222_ Shift_Register_Inst.data_out\[6\] Signal_Generator_1_90phase_inst.count\[1\]
+ _0241_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__and3b_1
X_1084_ _0493_ Dead_Time_Generator_inst_1.dt\[2\] net45 _0487_ VGND VGND VPWR VPWR
+ _0494_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0937_ _0403_ _0408_ net62 VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__a21oi_1
X_0799_ Signal_Generator_1_90phase_inst.count\[2\] _0298_ VGND VGND VPWR VPWR _0305_
+ sky130_fd_sc_hd__xor2_1
X_0868_ net77 _0355_ _0356_ _0340_ _0357_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0722_ _0215_ _0248_ _0223_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1136_ net9 _0538_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__and2b_1
X_1205_ _0242_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or2_1
X_1067_ _0485_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0705_ _0219_ _0220_ _0221_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__or3b_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1119_ _0525_ _0526_ _0522_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1470_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0193_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0970_ _0424_ _0431_ _0433_ Signal_Generator_2_270phase_inst.direction VGND VGND
+ VPWR VPWR _0052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1453_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0176_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[2\] sky130_fd_sc_hd__dfxtp_1
X_1384_ clknet_1_0__leaf_CLK_SR _0163_ _0084_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0953_ Signal_Generator_2_180phase_inst.count\[4\] Signal_Generator_2_180phase_inst.direction
+ _0401_ Signal_Generator_2_180phase_inst.count\[5\] VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__o31a_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0884_ Signal_Generator_2_0phase_inst.count\[2\] _0362_ VGND VGND VPWR VPWR _0369_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1436_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0062_ _0135_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_1367_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0000_ _0067_ VGND VGND VPWR
+ VPWR NMOS1_PS1_prev sky130_fd_sc_hd__dfrtp_1
X_1298_ _0633_ _0643_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1221_ Shift_Register_Inst.data_out\[5\] Shift_Register_Inst.data_out\[6\] Signal_Generator_1_180phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__and3b_1
Xclkbuf_1_1__f_CLK_SR clknet_0_CLK_SR VGND VGND VPWR VPWR clknet_1_1__leaf_CLK_SR
+ sky130_fd_sc_hd__clkbuf_16
X_1152_ _0551_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
X_1083_ Dead_Time_Generator_inst_4.count_dt\[2\] VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__inv_2
X_0936_ _0407_ _0404_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0798_ Signal_Generator_1_90phase_inst.count\[2\] _0301_ VGND VGND VPWR VPWR _0304_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0867_ Signal_Generator_1_270phase_inst.count\[4\] _0338_ VGND VGND VPWR VPWR _0357_
+ sky130_fd_sc_hd__xnor2_1
X_1419_ clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk _0024_ _0118_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[2\] sky130_fd_sc_hd__dfrtp_4
X_0721_ Shift_Register_Inst.data_out\[7\] VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__buf_2
X_1204_ Shift_Register_Inst.data_out\[6\] VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1135_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__buf_2
X_1066_ _0485_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
X_0919_ _0394_ _0395_ _0385_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 Shift_Register_Inst.data_out\[15\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0704_ _0235_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1049_ _0483_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__inv_2
X_1118_ _0519_ _0520_ _0515_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1452_ clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk _0175_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[1\] sky130_fd_sc_hd__dfxtp_1
X_1383_ clknet_1_0__leaf_CLK_SR _0162_ _0083_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0952_ net62 _0418_ _0419_ _0403_ _0420_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0883_ Signal_Generator_2_0phase_inst.count\[2\] _0365_ VGND VGND VPWR VPWR _0368_
+ sky130_fd_sc_hd__xor2_1
X_1435_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0061_ _0134_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[4\] sky130_fd_sc_hd__dfstp_2
X_1366_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk net32 _0066_ VGND VGND VPWR
+ VPWR PMOS2_PS1_prev sky130_fd_sc_hd__dfstp_1
X_1297_ Dead_Time_Generator_inst_2.count_dt\[0\] _0633_ _0643_ VGND VGND VPWR VPWR
+ _0644_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1151_ _0551_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
X_1220_ Signal_Generator_1_0phase_inst.count\[1\] _0558_ VGND VGND VPWR VPWR _0573_
+ sky130_fd_sc_hd__or2_1
X_1082_ _0488_ Dead_Time_Generator_inst_1.dt\[0\] _0489_ _0490_ _0491_ VGND VGND VPWR
+ VPWR _0492_ sky130_fd_sc_hd__a311o_1
X_0935_ Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__nor2_1
X_0866_ Signal_Generator_1_270phase_inst.count\[4\] _0342_ VGND VGND VPWR VPWR _0356_
+ sky130_fd_sc_hd__or2_1
X_0797_ _0035_ _0302_ _0303_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__a21oi_1
X_1349_ Dead_Time_Generator_inst_4.count_dt\[1\] _0201_ VGND VGND VPWR VPWR _0205_
+ sky130_fd_sc_hd__xor2_1
X_1418_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0023_ _0117_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0720_ _0247_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1203_ _0445_ net8 VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__nand2_1
X_1134_ _0511_ _0512_ _0514_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__a22o_1
X_1065_ _0482_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__buf_4
X_0918_ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__a31o_1
X_0849_ _0340_ _0343_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__nor2_1
Xhold6 net30 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
X_0703_ _0215_ Dead_Time_Generator_inst_1.dt\[2\] _0234_ VGND VGND VPWR VPWR _0235_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1117_ _0522_ _0525_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1048_ _0483_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1382_ clknet_1_1__leaf_CLK_SR _0161_ _0082_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_1451_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk net42 VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_1.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0951_ Signal_Generator_2_180phase_inst.count\[4\] _0401_ VGND VGND VPWR VPWR _0420_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0882_ _0042_ _0366_ _0367_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1434_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0060_ _0133_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[3\] sky130_fd_sc_hd__dfstp_1
X_1296_ _0634_ net39 _0639_ _0641_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a221o_1
X_1365_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0002_ _0065_ VGND VGND VPWR
+ VPWR NMOS2_PS1_prev sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ _0551_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
X_1081_ Dead_Time_Generator_inst_4.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0934_ net57 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
X_0865_ _0352_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__or3b_1
Xclkbuf_3_6__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
X_0796_ _0297_ _0302_ net63 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1417_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0022_ _0116_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.count\[0\] sky130_fd_sc_hd__dfrtp_2
X_1279_ _0614_ _0627_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1348_ _0204_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
X_1202_ _0482_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1064_ _0484_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
X_1133_ _0530_ _0541_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a21o_1
X_0917_ _0384_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__inv_2
X_0779_ _0276_ _0287_ _0290_ Signal_Generator_1_0phase_inst.direction VGND VGND VPWR
+ VPWR _0011_ sky130_fd_sc_hd__a22o_1
X_0848_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_CLK_SR CLK_SR VGND VGND VPWR VPWR clknet_0_CLK_SR sky130_fd_sc_hd__clkbuf_16
Xhold7 _0006_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
X_0702_ Shift_Register_Inst.shift_state\[3\] _0220_ _0233_ VGND VGND VPWR VPWR _0234_
+ sky130_fd_sc_hd__or3_1
X_1047_ _0483_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__inv_2
X_1116_ Signal_Generator_2_0phase_inst.count\[2\] _0498_ VGND VGND VPWR VPWR _0526_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1450_ clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk _0055_ _0149_ VGND VGND VPWR
+ VPWR Signal_Generator_2_270phase_inst.count\[5\] sky130_fd_sc_hd__dfstp_1
X_1381_ clknet_1_1__leaf_CLK_SR _0160_ _0081_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0950_ Signal_Generator_2_180phase_inst.count\[4\] _0405_ VGND VGND VPWR VPWR _0419_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0881_ _0361_ _0366_ net69 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__a21oi_1
X_1433_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0059_ _0132_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[2\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_10_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1295_ Dead_Time_Generator_inst_2.count_dt\[4\] net53 VGND VGND VPWR VPWR _0642_
+ sky130_fd_sc_hd__and2b_1
X_1364_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk net34 _0064_ VGND VGND VPWR
+ VPWR PMOS1_PS1_prev sky130_fd_sc_hd__dfstp_1
XFILLER_0_18_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1080_ Dead_Time_Generator_inst_4.count_dt\[2\] Dead_Time_Generator_inst_1.dt\[2\]
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__and2b_1
X_0933_ _0403_ _0406_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__nor2_1
X_0795_ _0301_ _0298_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or2_1
X_0864_ _0340_ _0351_ _0354_ net68 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1347_ _0545_ _0549_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__and3_1
X_1416_ clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk _0028_ _0115_ VGND VGND VPWR
+ VPWR Signal_Generator_1_270phase_inst.direction sky130_fd_sc_hd__dfrtp_1
X_1278_ _0625_ _0626_ _0629_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__a21oi_1
X_1201_ _0482_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1063_ _0484_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1132_ _0521_ _0527_ _0528_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__o21a_1
X_0916_ _0380_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__nand2_1
X_0778_ _0288_ _0289_ _0279_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a21o_1
X_0847_ Signal_Generator_1_270phase_inst.count\[3\] Signal_Generator_1_270phase_inst.count\[2\]
+ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold8 net85 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0701_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[0\]
+ Shift_Register_Inst.shift_state\[1\] VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or3b_1
XFILLER_0_45_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1115_ _0506_ Signal_Generator_2_90phase_inst.count\[2\] _0500_ _0523_ _0524_ VGND
+ VGND VPWR VPWR _0525_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1046_ _0483_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1029_ Dead_Time_Generator_inst_2.go net3 _0262_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1380_ clknet_1_0__leaf_CLK_SR _0159_ _0080_ VGND VGND VPWR VPWR Shift_Register_Inst.data_out\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0880_ _0365_ _0362_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__or2_1
X_1432_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0058_ _0131_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1363_ _0545_ _0549_ net38 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1294_ _0640_ Dead_Time_Generator_inst_1.dt\[2\] net45 _0634_ VGND VGND VPWR VPWR
+ _0641_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ Signal_Generator_2_180phase_inst.count\[5\] Signal_Generator_2_180phase_inst.count\[4\]
+ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0794_ Signal_Generator_1_90phase_inst.count\[0\] Signal_Generator_1_90phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nor2_1
X_0863_ _0352_ _0353_ _0343_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a21o_1
X_1346_ _0201_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__nor2_1
X_1415_ clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk _0020_ _0114_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[5\] sky130_fd_sc_hd__dfstp_1
X_1277_ _0627_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__nand2_1
X_1200_ _0482_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1062_ _0484_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_2
X_1131_ _0537_ _0539_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a21o_1
X_0915_ Signal_Generator_2_90phase_inst.count\[2\] Signal_Generator_2_90phase_inst.count\[1\]
+ Signal_Generator_2_90phase_inst.count\[0\] Signal_Generator_2_90phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_7_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0777_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a31o_1
X_0846_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__and2_1
X_1329_ _0659_ _0668_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__and2_1
Xhold9 _0004_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0700_ _0232_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_1114_ _0248_ _0250_ Signal_Generator_2_270phase_inst.count\[2\] VGND VGND VPWR VPWR
+ _0524_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1045_ _0483_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__inv_2
X_0829_ _0322_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1028_ net31 VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1431_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0057_ _0130_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_2
X_1293_ Dead_Time_Generator_inst_2.count_dt\[2\] VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1362_ _0214_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ Signal_Generator_2_180phase_inst.count\[3\] Signal_Generator_2_180phase_inst.count\[2\]
+ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__and3_1
X_0862_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[2\] Signal_Generator_1_270phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0793_ net60 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
X_1276_ Dead_Time_Generator_inst_1.count_dt\[1\] _0622_ VGND VGND VPWR VPWR _0628_
+ sky130_fd_sc_hd__or2_1
X_1414_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0019_ _0113_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[4\] sky130_fd_sc_hd__dfstp_2
X_1345_ _0488_ _0497_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1130_ _0536_ _0531_ _0535_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__and3_1
X_1061_ _0484_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
X_0914_ _0382_ _0389_ _0391_ net65 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a22o_1
X_0845_ Signal_Generator_1_270phase_inst.count\[5\] Signal_Generator_1_270phase_inst.count\[4\]
+ _0338_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o31a_1
X_0776_ _0278_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1259_ net37 Dead_Time_Generator_inst_1.count_dt\[4\] VGND VGND VPWR VPWR _0612_
+ sky130_fd_sc_hd__or2b_1
X_1328_ Dead_Time_Generator_inst_3.count_dt\[0\] _0659_ _0668_ VGND VGND VPWR VPWR
+ _0669_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ Shift_Register_Inst.data_out\[7\] _0250_ Signal_Generator_2_180phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__and3b_1
X_1044_ _0483_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0828_ Signal_Generator_1_180phase_inst.count\[2\] _0320_ VGND VGND VPWR VPWR _0327_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0759_ Signal_Generator_1_0phase_inst.direction VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1027_ _0262_ Dead_Time_Generator_inst_3.go _0473_ net31 VGND VGND VPWR VPWR _0006_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7__f_Dead_Time_Generator_inst_1.clk clknet_0_Dead_Time_Generator_inst_1.clk
+ VGND VGND VPWR VPWR clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1430_ clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk _0063_ _0129_ VGND VGND VPWR
+ VPWR Signal_Generator_2_90phase_inst.direction sky130_fd_sc_hd__dfstp_1
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1292_ _0635_ Dead_Time_Generator_inst_1.dt\[0\] _0636_ _0637_ _0638_ VGND VGND VPWR
+ VPWR _0639_ sky130_fd_sc_hd__a311o_1
X_1361_ _0545_ _0549_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0930_ Signal_Generator_2_180phase_inst.count\[1\] Signal_Generator_2_180phase_inst.count\[0\]
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__and2_1
X_0792_ _0297_ _0300_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__nor2_1
X_0861_ _0342_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__inv_2
X_1413_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0018_ _0112_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[3\] sky130_fd_sc_hd__dfstp_1
X_1275_ Dead_Time_Generator_inst_1.count_dt\[1\] _0622_ VGND VGND VPWR VPWR _0627_
+ sky130_fd_sc_hd__nand2_1
X_1344_ Dead_Time_Generator_inst_4.count_dt\[0\] _0486_ _0496_ VGND VGND VPWR VPWR
+ _0201_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1060_ _0484_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_2
X_0913_ _0385_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0775_ _0274_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nand2_1
X_0844_ Signal_Generator_1_270phase_inst.direction VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__inv_2
X_1189_ _0555_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1258_ _0608_ _0610_ _0601_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or3b_1
X_1327_ _0660_ net39 _0665_ _0666_ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1112_ net11 VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__inv_2
X_1043_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0827_ Signal_Generator_1_180phase_inst.count\[2\] _0323_ VGND VGND VPWR VPWR _0326_
+ sky130_fd_sc_hd__xor2_1
X_0758_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[3\] Signal_Generator_1_0phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__or4_2
X_0689_ _0220_ _0221_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1026_ _0262_ net4 VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ Shift_Register_Inst.data_out\[9\] Shift_Register_Inst.data_out\[10\] VGND
+ VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1360_ Dead_Time_Generator_inst_4.count_dt\[3\] _0207_ Dead_Time_Generator_inst_4.count_dt\[4\]
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1291_ Dead_Time_Generator_inst_2.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0791_ Signal_Generator_1_90phase_inst.count\[5\] Signal_Generator_1_90phase_inst.count\[4\]
+ _0299_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__and3_1
X_0860_ _0338_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__nand2_1
X_1412_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0017_ _0111_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[2\] sky130_fd_sc_hd__dfstp_2
X_1343_ _0200_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1274_ _0611_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__buf_2
X_0989_ _0446_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_0_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0912_ Signal_Generator_2_90phase_inst.count\[2\] _0383_ VGND VGND VPWR VPWR _0390_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0774_ Signal_Generator_1_0phase_inst.count\[0\] Signal_Generator_1_0phase_inst.count\[1\]
+ Signal_Generator_1_0phase_inst.count\[2\] Signal_Generator_1_0phase_inst.count\[3\]
+ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o31ai_1
X_0843_ Signal_Generator_1_270phase_inst.count\[0\] Signal_Generator_1_270phase_inst.count\[1\]
+ Signal_Generator_1_270phase_inst.count\[3\] Signal_Generator_1_270phase_inst.count\[2\]
+ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__or4_2
XFILLER_0_45_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1326_ Dead_Time_Generator_inst_3.count_dt\[4\] net37 VGND VGND VPWR VPWR _0667_
+ sky130_fd_sc_hd__and2b_1
X_1188_ _0555_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_2
X_1257_ _0563_ _0572_ _0605_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1111_ _0515_ _0519_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and3_1
X_1042_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0688_ _0223_ _0224_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__nand2_1
X_0757_ _0273_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0826_ _0021_ _0324_ _0325_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1309_ _0625_ _0626_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1025_ _0262_ Dead_Time_Generator_inst_1.go _0472_ net31 VGND VGND VPWR VPWR _0004_
+ sky130_fd_sc_hd__o211ai_1
X_0809_ _0312_ Signal_Generator_1_90phase_inst.count\[4\] _0299_ VGND VGND VPWR VPWR
+ _0313_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 CLK_EXT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ net19 _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1290_ Dead_Time_Generator_inst_2.count_dt\[2\] Dead_Time_Generator_inst_1.dt\[2\]
+ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0790_ Signal_Generator_1_90phase_inst.count\[3\] Signal_Generator_1_90phase_inst.count\[2\]
+ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1411_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0016_ _0110_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[1\] sky130_fd_sc_hd__dfstp_1
X_1342_ _0625_ _0626_ _0645_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__and3_1
X_1273_ _0607_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0988_ _0445_ net7 VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0911_ Signal_Generator_2_90phase_inst.count\[2\] _0386_ VGND VGND VPWR VPWR _0389_
+ sky130_fd_sc_hd__xor2_1
X_0842_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0321_ _0337_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0773_ _0276_ _0283_ _0285_ Signal_Generator_1_0phase_inst.direction VGND VGND VPWR
+ VPWR _0010_ sky130_fd_sc_hd__a22o_1
X_1256_ _0602_ _0587_ _0579_ _0586_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__or4bb_1
X_1325_ _0661_ Dead_Time_Generator_inst_1.dt\[2\] net39 _0660_ VGND VGND VPWR VPWR
+ _0666_ sky130_fd_sc_hd__o22a_1
X_1187_ _0555_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1110_ Signal_Generator_2_0phase_inst.count\[3\] _0498_ VGND VGND VPWR VPWR _0520_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1041_ net2 VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0825_ _0319_ _0324_ net66 VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0687_ _0219_ _0222_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__nand2_1
X_0756_ Shift_Register_Inst.data_out\[17\] net1 _0272_ VGND VGND VPWR VPWR _0273_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1308_ _0651_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__and2b_1
X_1239_ _0557_ Signal_Generator_1_90phase_inst.count\[3\] VGND VGND VPWR VPWR _0592_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1024_ _0262_ net6 VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__nand2_1
X_0808_ Signal_Generator_1_90phase_inst.count\[5\] VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__inv_2
X_0739_ net1 Shift_Register_Inst.data_out\[12\] _0260_ VGND VGND VPWR VPWR _0261_
+ sky130_fd_sc_hd__mux2_1
Xhold60 Shift_Register_Inst.data_out\[13\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 CLK_PLL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_CLK_SR clknet_0_CLK_SR VGND VGND VPWR VPWR clknet_1_0__leaf_CLK_SR
+ sky130_fd_sc_hd__clkbuf_16
X_1007_ Shift_Register_Inst.data_out\[10\] Shift_Register_Inst.data_out\[9\] VGND
+ VGND VPWR VPWR _0456_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1410_ clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk _0015_ _0109_ VGND VGND VPWR
+ VPWR Signal_Generator_1_180phase_inst.count\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1272_ _0607_ _0611_ _0622_ _0624_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a211oi_1
X_1341_ _0545_ _0549_ _0198_ net56 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__o2bb2a_1
X_0987_ net41 VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0910_ _0063_ _0387_ _0388_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a21oi_1
X_0841_ Signal_Generator_1_180phase_inst.count\[4\] Signal_Generator_1_180phase_inst.direction
+ _0317_ Signal_Generator_1_180phase_inst.count\[5\] VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o31a_1
X_0772_ _0279_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1186_ _0481_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__buf_4
X_1255_ _0583_ _0584_ _0585_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__and3_1
X_1324_ _0661_ Dead_Time_Generator_inst_1.dt\[2\] _0662_ _0663_ _0664_ VGND VGND VPWR
+ VPWR _0665_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1040_ _0262_ net35 _0473_ _0474_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0755_ Shift_Register_Inst.shift_state\[4\] Shift_Register_Inst.shift_state\[0\]
+ _0271_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__and3_1
X_0824_ _0323_ _0320_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0686_ _0219_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1307_ Dead_Time_Generator_inst_2.count_dt\[1\] _0644_ Dead_Time_Generator_inst_2.count_dt\[2\]
+ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__a21o_1
X_1238_ _0241_ _0557_ Signal_Generator_1_180phase_inst.count\[3\] VGND VGND VPWR VPWR
+ _0591_ sky130_fd_sc_hd__and3b_1
X_1169_ _0553_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1023_ _0457_ _0461_ _0465_ _0471_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__o211a_4
X_0807_ _0297_ _0308_ _0311_ net63 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0738_ _0259_ _0238_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold50 Signal_Generator_1_0phase_inst.direction VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 Dead_Time_Generator_inst_1.dt\[4\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ _0455_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ _0544_ _0548_ _0198_ _0199_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1271_ Dead_Time_Generator_inst_1.count_dt\[0\] _0623_ VGND VGND VPWR VPWR _0624_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0986_ _0444_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
X_1469_ clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk _0192_ VGND VGND VPWR VPWR
+ Dead_Time_Generator_inst_4.count_dt\[0\] sky130_fd_sc_hd__dfxtp_1
X_0840_ net82 _0334_ _0335_ _0319_ _0336_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a32o_1
X_0771_ Signal_Generator_1_0phase_inst.count\[2\] _0277_ VGND VGND VPWR VPWR _0284_
+ sky130_fd_sc_hd__xor2_1
X_1323_ Dead_Time_Generator_inst_3.count_dt\[1\] Dead_Time_Generator_inst_1.dt\[1\]
+ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and2b_1
X_1185_ _0554_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
X_1254_ _0564_ _0572_ _0604_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__a22o_1
X_0969_ _0427_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0685_ _0220_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__nand2_1
X_0823_ Signal_Generator_1_180phase_inst.count\[0\] Signal_Generator_1_180phase_inst.count\[1\]
+ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0754_ _0216_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__inv_2
X_1306_ Dead_Time_Generator_inst_2.count_dt\[2\] Dead_Time_Generator_inst_2.count_dt\[1\]
+ _0644_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__and3_1
X_1099_ Signal_Generator_2_180phase_inst.count\[5\] _0499_ _0500_ VGND VGND VPWR VPWR
+ _0509_ sky130_fd_sc_hd__a21o_1
X_1237_ _0241_ _0557_ Signal_Generator_1_270phase_inst.count\[3\] VGND VGND VPWR VPWR
+ _0590_ sky130_fd_sc_hd__and3_1
X_1168_ _0553_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ Shift_Register_Inst.data_out\[12\] _0470_ Shift_Register_Inst.data_out\[11\]
+ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__o21ai_1
X_0806_ _0309_ _0310_ _0300_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0737_ _0219_ _0220_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold40 Signal_Generator_2_90phase_inst.direction VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold51 Shift_Register_Inst.data_out\[14\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1005_ PMOS1_PS1_prev _0448_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

