// This is the unpowered netlist.
module Top (CLK_EXT,
    CLK_PLL,
    CLK_SR,
    Data_SR,
    NMOS1_PS1,
    NMOS1_PS2,
    NMOS2_PS1,
    NMOS2_PS2,
    NMOS_PS3,
    PMOS1_PS1,
    PMOS1_PS2,
    PMOS2_PS1,
    PMOS2_PS2,
    PMOS_PS3,
    RST,
    SIGNAL_OUTPUT,
    d1,
    d2);
 input CLK_EXT;
 input CLK_PLL;
 input CLK_SR;
 input Data_SR;
 output NMOS1_PS1;
 output NMOS1_PS2;
 output NMOS2_PS1;
 output NMOS2_PS2;
 output NMOS_PS3;
 output PMOS1_PS1;
 output PMOS1_PS2;
 output PMOS2_PS1;
 output PMOS2_PS2;
 output PMOS_PS3;
 input RST;
 output SIGNAL_OUTPUT;
 input [5:0] d1;
 input [5:0] d2;

 wire \Dead_Time_Generator_inst_1.clk ;
 wire \Dead_Time_Generator_inst_1.count_dt[0] ;
 wire \Dead_Time_Generator_inst_1.count_dt[1] ;
 wire \Dead_Time_Generator_inst_1.count_dt[2] ;
 wire \Dead_Time_Generator_inst_1.count_dt[3] ;
 wire \Dead_Time_Generator_inst_1.count_dt[4] ;
 wire \Dead_Time_Generator_inst_1.dt[0] ;
 wire \Dead_Time_Generator_inst_1.dt[1] ;
 wire \Dead_Time_Generator_inst_1.dt[2] ;
 wire \Dead_Time_Generator_inst_1.dt[3] ;
 wire \Dead_Time_Generator_inst_1.dt[4] ;
 wire \Dead_Time_Generator_inst_1.go ;
 wire \Dead_Time_Generator_inst_2.count_dt[0] ;
 wire \Dead_Time_Generator_inst_2.count_dt[1] ;
 wire \Dead_Time_Generator_inst_2.count_dt[2] ;
 wire \Dead_Time_Generator_inst_2.count_dt[3] ;
 wire \Dead_Time_Generator_inst_2.count_dt[4] ;
 wire \Dead_Time_Generator_inst_2.go ;
 wire \Dead_Time_Generator_inst_3.count_dt[0] ;
 wire \Dead_Time_Generator_inst_3.count_dt[1] ;
 wire \Dead_Time_Generator_inst_3.count_dt[2] ;
 wire \Dead_Time_Generator_inst_3.count_dt[3] ;
 wire \Dead_Time_Generator_inst_3.count_dt[4] ;
 wire \Dead_Time_Generator_inst_3.go ;
 wire \Dead_Time_Generator_inst_4.count_dt[0] ;
 wire \Dead_Time_Generator_inst_4.count_dt[1] ;
 wire \Dead_Time_Generator_inst_4.count_dt[2] ;
 wire \Dead_Time_Generator_inst_4.count_dt[3] ;
 wire \Dead_Time_Generator_inst_4.count_dt[4] ;
 wire \Dead_Time_Generator_inst_4.go ;
 wire NMOS1_PS1_prev;
 wire NMOS1_PS2_prev;
 wire NMOS2_PS1_prev;
 wire NMOS2_PS2_prev;
 wire PMOS1_PS1_prev;
 wire PMOS1_PS2_prev;
 wire PMOS2_PS1_prev;
 wire PMOS2_PS2_prev;
 wire \Shift_Register_Inst.data_out[10] ;
 wire \Shift_Register_Inst.data_out[11] ;
 wire \Shift_Register_Inst.data_out[12] ;
 wire \Shift_Register_Inst.data_out[13] ;
 wire \Shift_Register_Inst.data_out[14] ;
 wire \Shift_Register_Inst.data_out[15] ;
 wire \Shift_Register_Inst.data_out[16] ;
 wire \Shift_Register_Inst.data_out[17] ;
 wire \Shift_Register_Inst.data_out[5] ;
 wire \Shift_Register_Inst.data_out[6] ;
 wire \Shift_Register_Inst.data_out[7] ;
 wire \Shift_Register_Inst.data_out[8] ;
 wire \Shift_Register_Inst.data_out[9] ;
 wire \Shift_Register_Inst.shift_state[0] ;
 wire \Shift_Register_Inst.shift_state[1] ;
 wire \Shift_Register_Inst.shift_state[2] ;
 wire \Shift_Register_Inst.shift_state[3] ;
 wire \Shift_Register_Inst.shift_state[4] ;
 wire \Signal_Generator_1_0phase_inst.count[0] ;
 wire \Signal_Generator_1_0phase_inst.count[1] ;
 wire \Signal_Generator_1_0phase_inst.count[2] ;
 wire \Signal_Generator_1_0phase_inst.count[3] ;
 wire \Signal_Generator_1_0phase_inst.count[4] ;
 wire \Signal_Generator_1_0phase_inst.count[5] ;
 wire \Signal_Generator_1_0phase_inst.direction ;
 wire \Signal_Generator_1_180phase_inst.count[0] ;
 wire \Signal_Generator_1_180phase_inst.count[1] ;
 wire \Signal_Generator_1_180phase_inst.count[2] ;
 wire \Signal_Generator_1_180phase_inst.count[3] ;
 wire \Signal_Generator_1_180phase_inst.count[4] ;
 wire \Signal_Generator_1_180phase_inst.count[5] ;
 wire \Signal_Generator_1_180phase_inst.direction ;
 wire \Signal_Generator_1_270phase_inst.count[0] ;
 wire \Signal_Generator_1_270phase_inst.count[1] ;
 wire \Signal_Generator_1_270phase_inst.count[2] ;
 wire \Signal_Generator_1_270phase_inst.count[3] ;
 wire \Signal_Generator_1_270phase_inst.count[4] ;
 wire \Signal_Generator_1_270phase_inst.count[5] ;
 wire \Signal_Generator_1_270phase_inst.direction ;
 wire \Signal_Generator_1_90phase_inst.count[0] ;
 wire \Signal_Generator_1_90phase_inst.count[1] ;
 wire \Signal_Generator_1_90phase_inst.count[2] ;
 wire \Signal_Generator_1_90phase_inst.count[3] ;
 wire \Signal_Generator_1_90phase_inst.count[4] ;
 wire \Signal_Generator_1_90phase_inst.count[5] ;
 wire \Signal_Generator_1_90phase_inst.direction ;
 wire \Signal_Generator_2_0phase_inst.count[0] ;
 wire \Signal_Generator_2_0phase_inst.count[1] ;
 wire \Signal_Generator_2_0phase_inst.count[2] ;
 wire \Signal_Generator_2_0phase_inst.count[3] ;
 wire \Signal_Generator_2_0phase_inst.count[4] ;
 wire \Signal_Generator_2_0phase_inst.count[5] ;
 wire \Signal_Generator_2_0phase_inst.direction ;
 wire \Signal_Generator_2_180phase_inst.count[0] ;
 wire \Signal_Generator_2_180phase_inst.count[1] ;
 wire \Signal_Generator_2_180phase_inst.count[2] ;
 wire \Signal_Generator_2_180phase_inst.count[3] ;
 wire \Signal_Generator_2_180phase_inst.count[4] ;
 wire \Signal_Generator_2_180phase_inst.count[5] ;
 wire \Signal_Generator_2_180phase_inst.direction ;
 wire \Signal_Generator_2_270phase_inst.count[0] ;
 wire \Signal_Generator_2_270phase_inst.count[1] ;
 wire \Signal_Generator_2_270phase_inst.count[2] ;
 wire \Signal_Generator_2_270phase_inst.count[3] ;
 wire \Signal_Generator_2_270phase_inst.count[4] ;
 wire \Signal_Generator_2_270phase_inst.count[5] ;
 wire \Signal_Generator_2_270phase_inst.direction ;
 wire \Signal_Generator_2_90phase_inst.count[0] ;
 wire \Signal_Generator_2_90phase_inst.count[1] ;
 wire \Signal_Generator_2_90phase_inst.count[2] ;
 wire \Signal_Generator_2_90phase_inst.count[3] ;
 wire \Signal_Generator_2_90phase_inst.count[4] ;
 wire \Signal_Generator_2_90phase_inst.count[5] ;
 wire \Signal_Generator_2_90phase_inst.direction ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire clknet_0_CLK_SR;
 wire \clknet_0_Dead_Time_Generator_inst_1.clk ;
 wire clknet_1_0__leaf_CLK_SR;
 wire clknet_1_1__leaf_CLK_SR;
 wire \clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ;
 wire \clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ;
 wire \clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ;
 wire \clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ;
 wire \clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ;
 wire \clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ;
 wire \clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ;
 wire \clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(CLK_EXT));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(CLK_PLL));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__buf_2 _0676_ (.A(net1),
    .X(_0215_));
 sky130_fd_sc_hd__or3_2 _0677_ (.A(\Shift_Register_Inst.shift_state[3] ),
    .B(\Shift_Register_Inst.shift_state[2] ),
    .C(\Shift_Register_Inst.shift_state[1] ),
    .X(_0216_));
 sky130_fd_sc_hd__or3_1 _0678_ (.A(\Shift_Register_Inst.shift_state[4] ),
    .B(\Shift_Register_Inst.shift_state[0] ),
    .C(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0679_ (.A0(_0215_),
    .A1(\Dead_Time_Generator_inst_1.dt[0] ),
    .S(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_1 _0680_ (.A(_0218_),
    .X(_0179_));
 sky130_fd_sc_hd__buf_2 _0681_ (.A(\Shift_Register_Inst.shift_state[3] ),
    .X(_0219_));
 sky130_fd_sc_hd__buf_2 _0682_ (.A(\Shift_Register_Inst.shift_state[2] ),
    .X(_0220_));
 sky130_fd_sc_hd__a41o_1 _0683_ (.A1(_0219_),
    .A2(_0220_),
    .A3(\Shift_Register_Inst.shift_state[1] ),
    .A4(\Shift_Register_Inst.shift_state[0] ),
    .B1(net61),
    .X(_0172_));
 sky130_fd_sc_hd__and3b_1 _0684_ (.A_N(\Shift_Register_Inst.shift_state[4] ),
    .B(\Shift_Register_Inst.shift_state[1] ),
    .C(\Shift_Register_Inst.shift_state[0] ),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _0685_ (.A(_0220_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__or2_1 _0686_ (.A(_0219_),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _0687_ (.A(_0219_),
    .B(_0222_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _0688_ (.A(_0223_),
    .B(_0224_),
    .Y(_0171_));
 sky130_fd_sc_hd__or2_1 _0689_ (.A(_0220_),
    .B(_0221_),
    .X(_0225_));
 sky130_fd_sc_hd__and2_1 _0690_ (.A(_0222_),
    .B(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _0691_ (.A(_0226_),
    .X(_0170_));
 sky130_fd_sc_hd__inv_2 _0692_ (.A(\Shift_Register_Inst.shift_state[0] ),
    .Y(_0227_));
 sky130_fd_sc_hd__and2_1 _0693_ (.A(\Shift_Register_Inst.shift_state[4] ),
    .B(_0216_),
    .X(_0228_));
 sky130_fd_sc_hd__or3_2 _0694_ (.A(\Shift_Register_Inst.shift_state[1] ),
    .B(_0227_),
    .C(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__o21ai_1 _0695_ (.A1(net61),
    .A2(_0227_),
    .B1(net64),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _0696_ (.A(_0229_),
    .B(_0230_),
    .Y(_0169_));
 sky130_fd_sc_hd__xnor2_1 _0697_ (.A(net67),
    .B(_0228_),
    .Y(_0168_));
 sky130_fd_sc_hd__or3_1 _0698_ (.A(\Shift_Register_Inst.shift_state[4] ),
    .B(_0227_),
    .C(_0216_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(_0215_),
    .A1(\Dead_Time_Generator_inst_1.dt[1] ),
    .S(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_1 _0700_ (.A(_0232_),
    .X(_0167_));
 sky130_fd_sc_hd__or3b_1 _0701_ (.A(\Shift_Register_Inst.shift_state[4] ),
    .B(\Shift_Register_Inst.shift_state[0] ),
    .C_N(\Shift_Register_Inst.shift_state[1] ),
    .X(_0233_));
 sky130_fd_sc_hd__or3_1 _0702_ (.A(\Shift_Register_Inst.shift_state[3] ),
    .B(_0220_),
    .C(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0703_ (.A0(_0215_),
    .A1(\Dead_Time_Generator_inst_1.dt[2] ),
    .S(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__clkbuf_1 _0704_ (.A(_0235_),
    .X(_0166_));
 sky130_fd_sc_hd__or3b_1 _0705_ (.A(_0219_),
    .B(_0220_),
    .C_N(_0221_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _0706_ (.A0(_0215_),
    .A1(\Dead_Time_Generator_inst_1.dt[3] ),
    .S(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_1 _0707_ (.A(_0237_),
    .X(_0165_));
 sky130_fd_sc_hd__or3_1 _0708_ (.A(\Shift_Register_Inst.shift_state[1] ),
    .B(\Shift_Register_Inst.shift_state[0] ),
    .C(_0228_),
    .X(_0238_));
 sky130_fd_sc_hd__or3b_1 _0709_ (.A(_0238_),
    .B(_0219_),
    .C_N(\Shift_Register_Inst.shift_state[2] ),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(_0215_),
    .A1(\Dead_Time_Generator_inst_1.dt[4] ),
    .S(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _0711_ (.A(_0240_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_2 _0712_ (.A(\Shift_Register_Inst.data_out[5] ),
    .X(_0241_));
 sky130_fd_sc_hd__buf_2 _0713_ (.A(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__or3b_1 _0714_ (.A(_0229_),
    .B(_0219_),
    .C_N(\Shift_Register_Inst.shift_state[2] ),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0715_ (.A0(_0215_),
    .A1(_0242_),
    .S(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_1 _0716_ (.A(_0244_),
    .X(_0163_));
 sky130_fd_sc_hd__buf_2 _0717_ (.A(\Shift_Register_Inst.data_out[6] ),
    .X(_0245_));
 sky130_fd_sc_hd__or3b_1 _0718_ (.A(_0233_),
    .B(_0219_),
    .C_N(\Shift_Register_Inst.shift_state[2] ),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(_0215_),
    .A1(_0245_),
    .S(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _0720_ (.A(_0247_),
    .X(_0162_));
 sky130_fd_sc_hd__buf_2 _0721_ (.A(\Shift_Register_Inst.data_out[7] ),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _0722_ (.A0(_0215_),
    .A1(_0248_),
    .S(_0223_),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_1 _0723_ (.A(_0249_),
    .X(_0161_));
 sky130_fd_sc_hd__buf_2 _0724_ (.A(\Shift_Register_Inst.data_out[8] ),
    .X(_0250_));
 sky130_fd_sc_hd__or3b_1 _0725_ (.A(_0220_),
    .B(_0238_),
    .C_N(\Shift_Register_Inst.shift_state[3] ),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(_0215_),
    .A1(_0250_),
    .S(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_1 _0727_ (.A(_0252_),
    .X(_0160_));
 sky130_fd_sc_hd__or3b_1 _0728_ (.A(_0220_),
    .B(_0229_),
    .C_N(\Shift_Register_Inst.shift_state[3] ),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0729_ (.A0(_0215_),
    .A1(\Shift_Register_Inst.data_out[9] ),
    .S(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__clkbuf_1 _0730_ (.A(_0254_),
    .X(_0159_));
 sky130_fd_sc_hd__or3b_1 _0731_ (.A(\Shift_Register_Inst.shift_state[2] ),
    .B(_0233_),
    .C_N(\Shift_Register_Inst.shift_state[3] ),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(net1),
    .A1(\Shift_Register_Inst.data_out[10] ),
    .S(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__clkbuf_1 _0733_ (.A(_0256_),
    .X(_0158_));
 sky130_fd_sc_hd__and3b_1 _0734_ (.A_N(_0220_),
    .B(_0221_),
    .C(_0219_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(\Shift_Register_Inst.data_out[11] ),
    .A1(net1),
    .S(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__clkbuf_1 _0736_ (.A(_0258_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_1 _0737_ (.A(_0219_),
    .B(_0220_),
    .Y(_0259_));
 sky130_fd_sc_hd__or2_1 _0738_ (.A(_0259_),
    .B(_0238_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _0739_ (.A0(net1),
    .A1(\Shift_Register_Inst.data_out[12] ),
    .S(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__clkbuf_1 _0740_ (.A(_0261_),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_4 _0741_ (.A(net33),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _0742_ (.A(_0259_),
    .B(_0229_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(net1),
    .A1(_0262_),
    .S(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_1 _0744_ (.A(_0264_),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _0745_ (.A(_0259_),
    .B(_0233_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(net1),
    .A1(net76),
    .S(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0266_),
    .X(_0154_));
 sky130_fd_sc_hd__and3_1 _0748_ (.A(_0219_),
    .B(_0220_),
    .C(_0221_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _0749_ (.A0(net79),
    .A1(net1),
    .S(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_1 _0750_ (.A(_0268_),
    .X(_0153_));
 sky130_fd_sc_hd__or3b_1 _0751_ (.A(\Shift_Register_Inst.shift_state[0] ),
    .B(_0216_),
    .C_N(\Shift_Register_Inst.shift_state[4] ),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(net1),
    .A1(\Shift_Register_Inst.data_out[16] ),
    .S(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0270_),
    .X(_0152_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(_0216_),
    .Y(_0271_));
 sky130_fd_sc_hd__and3_1 _0755_ (.A(\Shift_Register_Inst.shift_state[4] ),
    .B(\Shift_Register_Inst.shift_state[0] ),
    .C(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(\Shift_Register_Inst.data_out[17] ),
    .A1(net1),
    .S(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0273_),
    .X(_0151_));
 sky130_fd_sc_hd__or4_2 _0758_ (.A(\Signal_Generator_1_0phase_inst.count[0] ),
    .B(\Signal_Generator_1_0phase_inst.count[1] ),
    .C(\Signal_Generator_1_0phase_inst.count[3] ),
    .D(\Signal_Generator_1_0phase_inst.count[2] ),
    .X(_0274_));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(\Signal_Generator_1_0phase_inst.direction ),
    .Y(_0275_));
 sky130_fd_sc_hd__o31a_1 _0760_ (.A1(\Signal_Generator_1_0phase_inst.count[5] ),
    .A2(\Signal_Generator_1_0phase_inst.count[4] ),
    .A3(_0274_),
    .B1(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _0761_ (.A(\Signal_Generator_1_0phase_inst.count[0] ),
    .B(\Signal_Generator_1_0phase_inst.count[1] ),
    .X(_0277_));
 sky130_fd_sc_hd__and3_1 _0762_ (.A(\Signal_Generator_1_0phase_inst.count[3] ),
    .B(\Signal_Generator_1_0phase_inst.count[2] ),
    .C(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__and3_1 _0763_ (.A(\Signal_Generator_1_0phase_inst.count[5] ),
    .B(\Signal_Generator_1_0phase_inst.count[4] ),
    .C(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_1 _0764_ (.A(_0276_),
    .B(_0279_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(net52),
    .Y(_0008_));
 sky130_fd_sc_hd__nor2_1 _0766_ (.A(\Signal_Generator_1_0phase_inst.count[0] ),
    .B(\Signal_Generator_1_0phase_inst.count[1] ),
    .Y(_0280_));
 sky130_fd_sc_hd__or2_1 _0767_ (.A(_0280_),
    .B(_0277_),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_1 _0768_ (.A1(_0276_),
    .A2(_0281_),
    .B1(net75),
    .Y(_0282_));
 sky130_fd_sc_hd__a21oi_1 _0769_ (.A1(_0014_),
    .A2(_0281_),
    .B1(_0282_),
    .Y(_0009_));
 sky130_fd_sc_hd__xor2_1 _0770_ (.A(\Signal_Generator_1_0phase_inst.count[2] ),
    .B(_0280_),
    .X(_0283_));
 sky130_fd_sc_hd__xor2_1 _0771_ (.A(\Signal_Generator_1_0phase_inst.count[2] ),
    .B(_0277_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _0772_ (.A(_0279_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__a22o_1 _0773_ (.A1(_0276_),
    .A2(_0283_),
    .B1(_0285_),
    .B2(\Signal_Generator_1_0phase_inst.direction ),
    .X(_0010_));
 sky130_fd_sc_hd__o31ai_1 _0774_ (.A1(\Signal_Generator_1_0phase_inst.count[0] ),
    .A2(\Signal_Generator_1_0phase_inst.count[1] ),
    .A3(\Signal_Generator_1_0phase_inst.count[2] ),
    .B1(\Signal_Generator_1_0phase_inst.count[3] ),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_1 _0775_ (.A(_0274_),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(_0278_),
    .Y(_0288_));
 sky130_fd_sc_hd__a31o_1 _0777_ (.A1(\Signal_Generator_1_0phase_inst.count[0] ),
    .A2(\Signal_Generator_1_0phase_inst.count[1] ),
    .A3(\Signal_Generator_1_0phase_inst.count[2] ),
    .B1(\Signal_Generator_1_0phase_inst.count[3] ),
    .X(_0289_));
 sky130_fd_sc_hd__a21o_1 _0778_ (.A1(_0288_),
    .A2(_0289_),
    .B1(_0279_),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_1 _0779_ (.A1(_0276_),
    .A2(_0287_),
    .B1(_0290_),
    .B2(\Signal_Generator_1_0phase_inst.direction ),
    .X(_0011_));
 sky130_fd_sc_hd__or3b_1 _0780_ (.A(_0288_),
    .B(\Signal_Generator_1_0phase_inst.count[5] ),
    .C_N(\Signal_Generator_1_0phase_inst.count[4] ),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _0781_ (.A(\Signal_Generator_1_0phase_inst.count[4] ),
    .B(_0278_),
    .X(_0292_));
 sky130_fd_sc_hd__xnor2_1 _0782_ (.A(\Signal_Generator_1_0phase_inst.count[4] ),
    .B(_0274_),
    .Y(_0293_));
 sky130_fd_sc_hd__a32o_1 _0783_ (.A1(\Signal_Generator_1_0phase_inst.direction ),
    .A2(_0291_),
    .A3(_0292_),
    .B1(_0276_),
    .B2(_0293_),
    .X(_0012_));
 sky130_fd_sc_hd__o31a_1 _0784_ (.A1(\Signal_Generator_1_0phase_inst.count[4] ),
    .A2(\Signal_Generator_1_0phase_inst.direction ),
    .A3(_0274_),
    .B1(\Signal_Generator_1_0phase_inst.count[5] ),
    .X(_0294_));
 sky130_fd_sc_hd__a31o_1 _0785_ (.A1(net73),
    .A2(\Signal_Generator_1_0phase_inst.direction ),
    .A3(_0278_),
    .B1(_0294_),
    .X(_0013_));
 sky130_fd_sc_hd__or4_2 _0786_ (.A(\Signal_Generator_1_90phase_inst.count[0] ),
    .B(\Signal_Generator_1_90phase_inst.count[1] ),
    .C(\Signal_Generator_1_90phase_inst.count[3] ),
    .D(\Signal_Generator_1_90phase_inst.count[2] ),
    .X(_0295_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(\Signal_Generator_1_90phase_inst.direction ),
    .Y(_0296_));
 sky130_fd_sc_hd__o31a_1 _0788_ (.A1(\Signal_Generator_1_90phase_inst.count[5] ),
    .A2(\Signal_Generator_1_90phase_inst.count[4] ),
    .A3(_0295_),
    .B1(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__and2_1 _0789_ (.A(\Signal_Generator_1_90phase_inst.count[0] ),
    .B(\Signal_Generator_1_90phase_inst.count[1] ),
    .X(_0298_));
 sky130_fd_sc_hd__and3_1 _0790_ (.A(\Signal_Generator_1_90phase_inst.count[3] ),
    .B(\Signal_Generator_1_90phase_inst.count[2] ),
    .C(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__and3_1 _0791_ (.A(\Signal_Generator_1_90phase_inst.count[5] ),
    .B(\Signal_Generator_1_90phase_inst.count[4] ),
    .C(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__nor2_1 _0792_ (.A(_0297_),
    .B(_0300_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(net60),
    .Y(_0029_));
 sky130_fd_sc_hd__nor2_1 _0794_ (.A(\Signal_Generator_1_90phase_inst.count[0] ),
    .B(\Signal_Generator_1_90phase_inst.count[1] ),
    .Y(_0301_));
 sky130_fd_sc_hd__or2_1 _0795_ (.A(_0301_),
    .B(_0298_),
    .X(_0302_));
 sky130_fd_sc_hd__a21oi_1 _0796_ (.A1(_0297_),
    .A2(_0302_),
    .B1(net63),
    .Y(_0303_));
 sky130_fd_sc_hd__a21oi_1 _0797_ (.A1(_0035_),
    .A2(_0302_),
    .B1(_0303_),
    .Y(_0030_));
 sky130_fd_sc_hd__xor2_1 _0798_ (.A(\Signal_Generator_1_90phase_inst.count[2] ),
    .B(_0301_),
    .X(_0304_));
 sky130_fd_sc_hd__xor2_1 _0799_ (.A(\Signal_Generator_1_90phase_inst.count[2] ),
    .B(_0298_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _0800_ (.A(_0300_),
    .B(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__a22o_1 _0801_ (.A1(_0297_),
    .A2(_0304_),
    .B1(_0306_),
    .B2(net63),
    .X(_0031_));
 sky130_fd_sc_hd__o31ai_1 _0802_ (.A1(\Signal_Generator_1_90phase_inst.count[0] ),
    .A2(\Signal_Generator_1_90phase_inst.count[1] ),
    .A3(\Signal_Generator_1_90phase_inst.count[2] ),
    .B1(\Signal_Generator_1_90phase_inst.count[3] ),
    .Y(_0307_));
 sky130_fd_sc_hd__nand2_1 _0803_ (.A(_0295_),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(_0299_),
    .Y(_0309_));
 sky130_fd_sc_hd__a31o_1 _0805_ (.A1(\Signal_Generator_1_90phase_inst.count[0] ),
    .A2(\Signal_Generator_1_90phase_inst.count[1] ),
    .A3(\Signal_Generator_1_90phase_inst.count[2] ),
    .B1(\Signal_Generator_1_90phase_inst.count[3] ),
    .X(_0310_));
 sky130_fd_sc_hd__a21o_1 _0806_ (.A1(_0309_),
    .A2(_0310_),
    .B1(_0300_),
    .X(_0311_));
 sky130_fd_sc_hd__a22o_1 _0807_ (.A1(_0297_),
    .A2(_0308_),
    .B1(_0311_),
    .B2(net63),
    .X(_0032_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(\Signal_Generator_1_90phase_inst.count[5] ),
    .Y(_0312_));
 sky130_fd_sc_hd__and3_1 _0809_ (.A(_0312_),
    .B(\Signal_Generator_1_90phase_inst.count[4] ),
    .C(_0299_),
    .X(_0313_));
 sky130_fd_sc_hd__o21ai_1 _0810_ (.A1(\Signal_Generator_1_90phase_inst.count[4] ),
    .A2(_0299_),
    .B1(\Signal_Generator_1_90phase_inst.direction ),
    .Y(_0314_));
 sky130_fd_sc_hd__xnor2_1 _0811_ (.A(\Signal_Generator_1_90phase_inst.count[4] ),
    .B(_0295_),
    .Y(_0315_));
 sky130_fd_sc_hd__a2bb2o_1 _0812_ (.A1_N(_0313_),
    .A2_N(_0314_),
    .B1(_0297_),
    .B2(_0315_),
    .X(_0033_));
 sky130_fd_sc_hd__o31a_1 _0813_ (.A1(\Signal_Generator_1_90phase_inst.count[4] ),
    .A2(\Signal_Generator_1_90phase_inst.direction ),
    .A3(_0295_),
    .B1(\Signal_Generator_1_90phase_inst.count[5] ),
    .X(_0316_));
 sky130_fd_sc_hd__a31o_1 _0814_ (.A1(\Signal_Generator_1_90phase_inst.count[4] ),
    .A2(\Signal_Generator_1_90phase_inst.direction ),
    .A3(_0299_),
    .B1(_0316_),
    .X(_0034_));
 sky130_fd_sc_hd__or4_2 _0815_ (.A(\Signal_Generator_1_180phase_inst.count[0] ),
    .B(\Signal_Generator_1_180phase_inst.count[1] ),
    .C(\Signal_Generator_1_180phase_inst.count[3] ),
    .D(\Signal_Generator_1_180phase_inst.count[2] ),
    .X(_0317_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(\Signal_Generator_1_180phase_inst.direction ),
    .Y(_0318_));
 sky130_fd_sc_hd__o31a_2 _0817_ (.A1(\Signal_Generator_1_180phase_inst.count[5] ),
    .A2(\Signal_Generator_1_180phase_inst.count[4] ),
    .A3(_0317_),
    .B1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__and2_1 _0818_ (.A(\Signal_Generator_1_180phase_inst.count[0] ),
    .B(\Signal_Generator_1_180phase_inst.count[1] ),
    .X(_0320_));
 sky130_fd_sc_hd__and3_1 _0819_ (.A(\Signal_Generator_1_180phase_inst.count[3] ),
    .B(\Signal_Generator_1_180phase_inst.count[2] ),
    .C(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__and3_1 _0820_ (.A(\Signal_Generator_1_180phase_inst.count[5] ),
    .B(\Signal_Generator_1_180phase_inst.count[4] ),
    .C(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_1 _0821_ (.A(_0319_),
    .B(_0322_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(net59),
    .Y(_0015_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(\Signal_Generator_1_180phase_inst.count[0] ),
    .B(\Signal_Generator_1_180phase_inst.count[1] ),
    .Y(_0323_));
 sky130_fd_sc_hd__or2_1 _0824_ (.A(_0323_),
    .B(_0320_),
    .X(_0324_));
 sky130_fd_sc_hd__a21oi_1 _0825_ (.A1(_0319_),
    .A2(_0324_),
    .B1(net66),
    .Y(_0325_));
 sky130_fd_sc_hd__a21oi_1 _0826_ (.A1(_0021_),
    .A2(_0324_),
    .B1(_0325_),
    .Y(_0016_));
 sky130_fd_sc_hd__xor2_1 _0827_ (.A(\Signal_Generator_1_180phase_inst.count[2] ),
    .B(_0323_),
    .X(_0326_));
 sky130_fd_sc_hd__xor2_1 _0828_ (.A(\Signal_Generator_1_180phase_inst.count[2] ),
    .B(_0320_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _0829_ (.A(_0322_),
    .B(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _0830_ (.A1(_0319_),
    .A2(_0326_),
    .B1(_0328_),
    .B2(net66),
    .X(_0017_));
 sky130_fd_sc_hd__o31ai_1 _0831_ (.A1(\Signal_Generator_1_180phase_inst.count[0] ),
    .A2(\Signal_Generator_1_180phase_inst.count[1] ),
    .A3(\Signal_Generator_1_180phase_inst.count[2] ),
    .B1(\Signal_Generator_1_180phase_inst.count[3] ),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_1 _0832_ (.A(_0317_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(_0321_),
    .Y(_0331_));
 sky130_fd_sc_hd__a31o_1 _0834_ (.A1(\Signal_Generator_1_180phase_inst.count[0] ),
    .A2(\Signal_Generator_1_180phase_inst.count[1] ),
    .A3(\Signal_Generator_1_180phase_inst.count[2] ),
    .B1(\Signal_Generator_1_180phase_inst.count[3] ),
    .X(_0332_));
 sky130_fd_sc_hd__a21o_1 _0835_ (.A1(_0331_),
    .A2(_0332_),
    .B1(_0322_),
    .X(_0333_));
 sky130_fd_sc_hd__a22o_1 _0836_ (.A1(_0319_),
    .A2(_0330_),
    .B1(_0333_),
    .B2(net66),
    .X(_0018_));
 sky130_fd_sc_hd__or3b_1 _0837_ (.A(_0331_),
    .B(\Signal_Generator_1_180phase_inst.count[5] ),
    .C_N(\Signal_Generator_1_180phase_inst.count[4] ),
    .X(_0334_));
 sky130_fd_sc_hd__or2_1 _0838_ (.A(\Signal_Generator_1_180phase_inst.count[4] ),
    .B(_0321_),
    .X(_0335_));
 sky130_fd_sc_hd__xnor2_1 _0839_ (.A(\Signal_Generator_1_180phase_inst.count[4] ),
    .B(_0317_),
    .Y(_0336_));
 sky130_fd_sc_hd__a32o_1 _0840_ (.A1(net82),
    .A2(_0334_),
    .A3(_0335_),
    .B1(_0319_),
    .B2(_0336_),
    .X(_0019_));
 sky130_fd_sc_hd__o31a_1 _0841_ (.A1(\Signal_Generator_1_180phase_inst.count[4] ),
    .A2(\Signal_Generator_1_180phase_inst.direction ),
    .A3(_0317_),
    .B1(\Signal_Generator_1_180phase_inst.count[5] ),
    .X(_0337_));
 sky130_fd_sc_hd__a31o_1 _0842_ (.A1(\Signal_Generator_1_180phase_inst.count[4] ),
    .A2(\Signal_Generator_1_180phase_inst.direction ),
    .A3(_0321_),
    .B1(_0337_),
    .X(_0020_));
 sky130_fd_sc_hd__or4_2 _0843_ (.A(\Signal_Generator_1_270phase_inst.count[0] ),
    .B(\Signal_Generator_1_270phase_inst.count[1] ),
    .C(\Signal_Generator_1_270phase_inst.count[3] ),
    .D(\Signal_Generator_1_270phase_inst.count[2] ),
    .X(_0338_));
 sky130_fd_sc_hd__inv_2 _0844_ (.A(\Signal_Generator_1_270phase_inst.direction ),
    .Y(_0339_));
 sky130_fd_sc_hd__o31a_1 _0845_ (.A1(\Signal_Generator_1_270phase_inst.count[5] ),
    .A2(\Signal_Generator_1_270phase_inst.count[4] ),
    .A3(_0338_),
    .B1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__and2_1 _0846_ (.A(\Signal_Generator_1_270phase_inst.count[0] ),
    .B(\Signal_Generator_1_270phase_inst.count[1] ),
    .X(_0341_));
 sky130_fd_sc_hd__and3_1 _0847_ (.A(\Signal_Generator_1_270phase_inst.count[3] ),
    .B(\Signal_Generator_1_270phase_inst.count[2] ),
    .C(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__and3_1 _0848_ (.A(\Signal_Generator_1_270phase_inst.count[5] ),
    .B(\Signal_Generator_1_270phase_inst.count[4] ),
    .C(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__nor2_1 _0849_ (.A(_0340_),
    .B(_0343_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0850_ (.A(net48),
    .Y(_0022_));
 sky130_fd_sc_hd__nor2_1 _0851_ (.A(\Signal_Generator_1_270phase_inst.count[0] ),
    .B(\Signal_Generator_1_270phase_inst.count[1] ),
    .Y(_0344_));
 sky130_fd_sc_hd__or2_1 _0852_ (.A(_0344_),
    .B(_0341_),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_1 _0853_ (.A1(_0340_),
    .A2(_0345_),
    .B1(net68),
    .Y(_0346_));
 sky130_fd_sc_hd__a21oi_1 _0854_ (.A1(_0028_),
    .A2(_0345_),
    .B1(_0346_),
    .Y(_0023_));
 sky130_fd_sc_hd__xor2_1 _0855_ (.A(\Signal_Generator_1_270phase_inst.count[2] ),
    .B(_0344_),
    .X(_0347_));
 sky130_fd_sc_hd__xor2_1 _0856_ (.A(\Signal_Generator_1_270phase_inst.count[2] ),
    .B(_0341_),
    .X(_0348_));
 sky130_fd_sc_hd__or2_1 _0857_ (.A(_0343_),
    .B(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__a22o_1 _0858_ (.A1(_0340_),
    .A2(_0347_),
    .B1(_0349_),
    .B2(net68),
    .X(_0024_));
 sky130_fd_sc_hd__o31ai_1 _0859_ (.A1(\Signal_Generator_1_270phase_inst.count[0] ),
    .A2(\Signal_Generator_1_270phase_inst.count[1] ),
    .A3(\Signal_Generator_1_270phase_inst.count[2] ),
    .B1(\Signal_Generator_1_270phase_inst.count[3] ),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _0860_ (.A(_0338_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _0861_ (.A(_0342_),
    .Y(_0352_));
 sky130_fd_sc_hd__a31o_1 _0862_ (.A1(\Signal_Generator_1_270phase_inst.count[0] ),
    .A2(\Signal_Generator_1_270phase_inst.count[1] ),
    .A3(\Signal_Generator_1_270phase_inst.count[2] ),
    .B1(\Signal_Generator_1_270phase_inst.count[3] ),
    .X(_0353_));
 sky130_fd_sc_hd__a21o_1 _0863_ (.A1(_0352_),
    .A2(_0353_),
    .B1(_0343_),
    .X(_0354_));
 sky130_fd_sc_hd__a22o_1 _0864_ (.A1(_0340_),
    .A2(_0351_),
    .B1(_0354_),
    .B2(net68),
    .X(_0025_));
 sky130_fd_sc_hd__or3b_1 _0865_ (.A(_0352_),
    .B(\Signal_Generator_1_270phase_inst.count[5] ),
    .C_N(\Signal_Generator_1_270phase_inst.count[4] ),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _0866_ (.A(\Signal_Generator_1_270phase_inst.count[4] ),
    .B(_0342_),
    .X(_0356_));
 sky130_fd_sc_hd__xnor2_1 _0867_ (.A(\Signal_Generator_1_270phase_inst.count[4] ),
    .B(_0338_),
    .Y(_0357_));
 sky130_fd_sc_hd__a32o_1 _0868_ (.A1(net77),
    .A2(_0355_),
    .A3(_0356_),
    .B1(_0340_),
    .B2(_0357_),
    .X(_0026_));
 sky130_fd_sc_hd__o31a_1 _0869_ (.A1(\Signal_Generator_1_270phase_inst.count[4] ),
    .A2(\Signal_Generator_1_270phase_inst.direction ),
    .A3(_0338_),
    .B1(\Signal_Generator_1_270phase_inst.count[5] ),
    .X(_0358_));
 sky130_fd_sc_hd__a31o_1 _0870_ (.A1(\Signal_Generator_1_270phase_inst.count[4] ),
    .A2(net77),
    .A3(_0342_),
    .B1(_0358_),
    .X(_0027_));
 sky130_fd_sc_hd__or4_2 _0871_ (.A(\Signal_Generator_2_0phase_inst.count[3] ),
    .B(\Signal_Generator_2_0phase_inst.count[2] ),
    .C(\Signal_Generator_2_0phase_inst.count[1] ),
    .D(\Signal_Generator_2_0phase_inst.count[0] ),
    .X(_0359_));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(\Signal_Generator_2_0phase_inst.direction ),
    .Y(_0360_));
 sky130_fd_sc_hd__o31a_1 _0873_ (.A1(\Signal_Generator_2_0phase_inst.count[5] ),
    .A2(\Signal_Generator_2_0phase_inst.count[4] ),
    .A3(_0359_),
    .B1(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _0874_ (.A(\Signal_Generator_2_0phase_inst.count[1] ),
    .B(\Signal_Generator_2_0phase_inst.count[0] ),
    .X(_0362_));
 sky130_fd_sc_hd__and3_1 _0875_ (.A(\Signal_Generator_2_0phase_inst.count[3] ),
    .B(\Signal_Generator_2_0phase_inst.count[2] ),
    .C(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__and3_1 _0876_ (.A(\Signal_Generator_2_0phase_inst.count[5] ),
    .B(\Signal_Generator_2_0phase_inst.count[4] ),
    .C(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__nor2_1 _0877_ (.A(_0361_),
    .B(_0364_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0878_ (.A(net58),
    .Y(_0036_));
 sky130_fd_sc_hd__nor2_1 _0879_ (.A(\Signal_Generator_2_0phase_inst.count[1] ),
    .B(\Signal_Generator_2_0phase_inst.count[0] ),
    .Y(_0365_));
 sky130_fd_sc_hd__or2_1 _0880_ (.A(_0365_),
    .B(_0362_),
    .X(_0366_));
 sky130_fd_sc_hd__a21oi_1 _0881_ (.A1(_0361_),
    .A2(_0366_),
    .B1(net69),
    .Y(_0367_));
 sky130_fd_sc_hd__a21oi_1 _0882_ (.A1(_0042_),
    .A2(_0366_),
    .B1(_0367_),
    .Y(_0037_));
 sky130_fd_sc_hd__xor2_1 _0883_ (.A(\Signal_Generator_2_0phase_inst.count[2] ),
    .B(_0365_),
    .X(_0368_));
 sky130_fd_sc_hd__xor2_1 _0884_ (.A(\Signal_Generator_2_0phase_inst.count[2] ),
    .B(_0362_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _0885_ (.A(_0364_),
    .B(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _0886_ (.A1(_0361_),
    .A2(_0368_),
    .B1(_0370_),
    .B2(net69),
    .X(_0038_));
 sky130_fd_sc_hd__o31ai_1 _0887_ (.A1(\Signal_Generator_2_0phase_inst.count[2] ),
    .A2(\Signal_Generator_2_0phase_inst.count[1] ),
    .A3(\Signal_Generator_2_0phase_inst.count[0] ),
    .B1(\Signal_Generator_2_0phase_inst.count[3] ),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _0888_ (.A(_0359_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _0889_ (.A(_0363_),
    .Y(_0373_));
 sky130_fd_sc_hd__a31o_1 _0890_ (.A1(\Signal_Generator_2_0phase_inst.count[2] ),
    .A2(\Signal_Generator_2_0phase_inst.count[1] ),
    .A3(\Signal_Generator_2_0phase_inst.count[0] ),
    .B1(\Signal_Generator_2_0phase_inst.count[3] ),
    .X(_0374_));
 sky130_fd_sc_hd__a21o_1 _0891_ (.A1(_0373_),
    .A2(_0374_),
    .B1(_0364_),
    .X(_0375_));
 sky130_fd_sc_hd__a22o_1 _0892_ (.A1(_0361_),
    .A2(_0372_),
    .B1(_0375_),
    .B2(net80),
    .X(_0039_));
 sky130_fd_sc_hd__or3b_1 _0893_ (.A(_0373_),
    .B(\Signal_Generator_2_0phase_inst.count[5] ),
    .C_N(\Signal_Generator_2_0phase_inst.count[4] ),
    .X(_0376_));
 sky130_fd_sc_hd__or2_1 _0894_ (.A(\Signal_Generator_2_0phase_inst.count[4] ),
    .B(_0363_),
    .X(_0377_));
 sky130_fd_sc_hd__xnor2_1 _0895_ (.A(\Signal_Generator_2_0phase_inst.count[4] ),
    .B(_0359_),
    .Y(_0378_));
 sky130_fd_sc_hd__a32o_1 _0896_ (.A1(net69),
    .A2(_0376_),
    .A3(_0377_),
    .B1(_0361_),
    .B2(_0378_),
    .X(_0040_));
 sky130_fd_sc_hd__o31a_1 _0897_ (.A1(\Signal_Generator_2_0phase_inst.count[4] ),
    .A2(\Signal_Generator_2_0phase_inst.direction ),
    .A3(_0359_),
    .B1(\Signal_Generator_2_0phase_inst.count[5] ),
    .X(_0379_));
 sky130_fd_sc_hd__a31o_1 _0898_ (.A1(\Signal_Generator_2_0phase_inst.count[4] ),
    .A2(\Signal_Generator_2_0phase_inst.direction ),
    .A3(_0363_),
    .B1(_0379_),
    .X(_0041_));
 sky130_fd_sc_hd__or4_2 _0899_ (.A(\Signal_Generator_2_90phase_inst.count[3] ),
    .B(\Signal_Generator_2_90phase_inst.count[2] ),
    .C(\Signal_Generator_2_90phase_inst.count[1] ),
    .D(\Signal_Generator_2_90phase_inst.count[0] ),
    .X(_0380_));
 sky130_fd_sc_hd__inv_2 _0900_ (.A(\Signal_Generator_2_90phase_inst.direction ),
    .Y(_0381_));
 sky130_fd_sc_hd__o31a_1 _0901_ (.A1(\Signal_Generator_2_90phase_inst.count[5] ),
    .A2(\Signal_Generator_2_90phase_inst.count[4] ),
    .A3(_0380_),
    .B1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _0902_ (.A(\Signal_Generator_2_90phase_inst.count[1] ),
    .B(\Signal_Generator_2_90phase_inst.count[0] ),
    .X(_0383_));
 sky130_fd_sc_hd__and3_1 _0903_ (.A(\Signal_Generator_2_90phase_inst.count[3] ),
    .B(\Signal_Generator_2_90phase_inst.count[2] ),
    .C(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__and3_1 _0904_ (.A(\Signal_Generator_2_90phase_inst.count[5] ),
    .B(\Signal_Generator_2_90phase_inst.count[4] ),
    .C(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_1 _0905_ (.A(_0382_),
    .B(_0385_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _0906_ (.A(net51),
    .Y(_0057_));
 sky130_fd_sc_hd__nor2_1 _0907_ (.A(\Signal_Generator_2_90phase_inst.count[1] ),
    .B(\Signal_Generator_2_90phase_inst.count[0] ),
    .Y(_0386_));
 sky130_fd_sc_hd__or2_1 _0908_ (.A(_0386_),
    .B(_0383_),
    .X(_0387_));
 sky130_fd_sc_hd__a21oi_1 _0909_ (.A1(_0382_),
    .A2(_0387_),
    .B1(net65),
    .Y(_0388_));
 sky130_fd_sc_hd__a21oi_1 _0910_ (.A1(_0063_),
    .A2(_0387_),
    .B1(_0388_),
    .Y(_0058_));
 sky130_fd_sc_hd__xor2_1 _0911_ (.A(\Signal_Generator_2_90phase_inst.count[2] ),
    .B(_0386_),
    .X(_0389_));
 sky130_fd_sc_hd__xor2_1 _0912_ (.A(\Signal_Generator_2_90phase_inst.count[2] ),
    .B(_0383_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _0913_ (.A(_0385_),
    .B(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(_0382_),
    .A2(_0389_),
    .B1(_0391_),
    .B2(net65),
    .X(_0059_));
 sky130_fd_sc_hd__o31ai_1 _0915_ (.A1(\Signal_Generator_2_90phase_inst.count[2] ),
    .A2(\Signal_Generator_2_90phase_inst.count[1] ),
    .A3(\Signal_Generator_2_90phase_inst.count[0] ),
    .B1(\Signal_Generator_2_90phase_inst.count[3] ),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _0916_ (.A(_0380_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__inv_2 _0917_ (.A(_0384_),
    .Y(_0394_));
 sky130_fd_sc_hd__a31o_1 _0918_ (.A1(\Signal_Generator_2_90phase_inst.count[2] ),
    .A2(\Signal_Generator_2_90phase_inst.count[1] ),
    .A3(\Signal_Generator_2_90phase_inst.count[0] ),
    .B1(\Signal_Generator_2_90phase_inst.count[3] ),
    .X(_0395_));
 sky130_fd_sc_hd__a21o_1 _0919_ (.A1(_0394_),
    .A2(_0395_),
    .B1(_0385_),
    .X(_0396_));
 sky130_fd_sc_hd__a22o_1 _0920_ (.A1(_0382_),
    .A2(_0393_),
    .B1(_0396_),
    .B2(net65),
    .X(_0060_));
 sky130_fd_sc_hd__or3b_1 _0921_ (.A(_0394_),
    .B(\Signal_Generator_2_90phase_inst.count[5] ),
    .C_N(\Signal_Generator_2_90phase_inst.count[4] ),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _0922_ (.A(\Signal_Generator_2_90phase_inst.count[4] ),
    .B(_0384_),
    .X(_0398_));
 sky130_fd_sc_hd__xnor2_1 _0923_ (.A(\Signal_Generator_2_90phase_inst.count[4] ),
    .B(_0380_),
    .Y(_0399_));
 sky130_fd_sc_hd__a32o_1 _0924_ (.A1(net81),
    .A2(_0397_),
    .A3(_0398_),
    .B1(_0382_),
    .B2(_0399_),
    .X(_0061_));
 sky130_fd_sc_hd__o31a_1 _0925_ (.A1(\Signal_Generator_2_90phase_inst.count[4] ),
    .A2(\Signal_Generator_2_90phase_inst.direction ),
    .A3(_0380_),
    .B1(\Signal_Generator_2_90phase_inst.count[5] ),
    .X(_0400_));
 sky130_fd_sc_hd__a31o_1 _0926_ (.A1(\Signal_Generator_2_90phase_inst.count[4] ),
    .A2(\Signal_Generator_2_90phase_inst.direction ),
    .A3(_0384_),
    .B1(_0400_),
    .X(_0062_));
 sky130_fd_sc_hd__or4_2 _0927_ (.A(\Signal_Generator_2_180phase_inst.count[3] ),
    .B(\Signal_Generator_2_180phase_inst.count[2] ),
    .C(\Signal_Generator_2_180phase_inst.count[1] ),
    .D(\Signal_Generator_2_180phase_inst.count[0] ),
    .X(_0401_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(\Signal_Generator_2_180phase_inst.direction ),
    .Y(_0402_));
 sky130_fd_sc_hd__o31a_2 _0929_ (.A1(\Signal_Generator_2_180phase_inst.count[5] ),
    .A2(\Signal_Generator_2_180phase_inst.count[4] ),
    .A3(_0401_),
    .B1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__and2_1 _0930_ (.A(\Signal_Generator_2_180phase_inst.count[1] ),
    .B(\Signal_Generator_2_180phase_inst.count[0] ),
    .X(_0404_));
 sky130_fd_sc_hd__and3_1 _0931_ (.A(\Signal_Generator_2_180phase_inst.count[3] ),
    .B(\Signal_Generator_2_180phase_inst.count[2] ),
    .C(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__and3_1 _0932_ (.A(\Signal_Generator_2_180phase_inst.count[5] ),
    .B(\Signal_Generator_2_180phase_inst.count[4] ),
    .C(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_1 _0933_ (.A(_0403_),
    .B(_0406_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(net57),
    .Y(_0043_));
 sky130_fd_sc_hd__nor2_1 _0935_ (.A(\Signal_Generator_2_180phase_inst.count[1] ),
    .B(\Signal_Generator_2_180phase_inst.count[0] ),
    .Y(_0407_));
 sky130_fd_sc_hd__or2_1 _0936_ (.A(_0407_),
    .B(_0404_),
    .X(_0408_));
 sky130_fd_sc_hd__a21oi_1 _0937_ (.A1(_0403_),
    .A2(_0408_),
    .B1(net62),
    .Y(_0409_));
 sky130_fd_sc_hd__a21oi_1 _0938_ (.A1(_0049_),
    .A2(_0408_),
    .B1(_0409_),
    .Y(_0044_));
 sky130_fd_sc_hd__xor2_1 _0939_ (.A(\Signal_Generator_2_180phase_inst.count[2] ),
    .B(_0407_),
    .X(_0410_));
 sky130_fd_sc_hd__xor2_1 _0940_ (.A(\Signal_Generator_2_180phase_inst.count[2] ),
    .B(_0404_),
    .X(_0411_));
 sky130_fd_sc_hd__or2_1 _0941_ (.A(_0406_),
    .B(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _0942_ (.A1(_0403_),
    .A2(_0410_),
    .B1(_0412_),
    .B2(net62),
    .X(_0045_));
 sky130_fd_sc_hd__o31ai_1 _0943_ (.A1(\Signal_Generator_2_180phase_inst.count[2] ),
    .A2(\Signal_Generator_2_180phase_inst.count[1] ),
    .A3(\Signal_Generator_2_180phase_inst.count[0] ),
    .B1(\Signal_Generator_2_180phase_inst.count[3] ),
    .Y(_0413_));
 sky130_fd_sc_hd__nand2_1 _0944_ (.A(_0401_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_2 _0945_ (.A(_0405_),
    .Y(_0415_));
 sky130_fd_sc_hd__a31o_1 _0946_ (.A1(\Signal_Generator_2_180phase_inst.count[2] ),
    .A2(\Signal_Generator_2_180phase_inst.count[1] ),
    .A3(\Signal_Generator_2_180phase_inst.count[0] ),
    .B1(\Signal_Generator_2_180phase_inst.count[3] ),
    .X(_0416_));
 sky130_fd_sc_hd__a21o_1 _0947_ (.A1(_0415_),
    .A2(_0416_),
    .B1(_0406_),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _0948_ (.A1(_0403_),
    .A2(_0414_),
    .B1(_0417_),
    .B2(net62),
    .X(_0046_));
 sky130_fd_sc_hd__or3b_1 _0949_ (.A(_0415_),
    .B(\Signal_Generator_2_180phase_inst.count[5] ),
    .C_N(\Signal_Generator_2_180phase_inst.count[4] ),
    .X(_0418_));
 sky130_fd_sc_hd__or2_1 _0950_ (.A(\Signal_Generator_2_180phase_inst.count[4] ),
    .B(_0405_),
    .X(_0419_));
 sky130_fd_sc_hd__xnor2_1 _0951_ (.A(\Signal_Generator_2_180phase_inst.count[4] ),
    .B(_0401_),
    .Y(_0420_));
 sky130_fd_sc_hd__a32o_1 _0952_ (.A1(net62),
    .A2(_0418_),
    .A3(_0419_),
    .B1(_0403_),
    .B2(_0420_),
    .X(_0047_));
 sky130_fd_sc_hd__o31a_1 _0953_ (.A1(\Signal_Generator_2_180phase_inst.count[4] ),
    .A2(\Signal_Generator_2_180phase_inst.direction ),
    .A3(_0401_),
    .B1(\Signal_Generator_2_180phase_inst.count[5] ),
    .X(_0421_));
 sky130_fd_sc_hd__a31o_1 _0954_ (.A1(\Signal_Generator_2_180phase_inst.count[4] ),
    .A2(net83),
    .A3(_0405_),
    .B1(_0421_),
    .X(_0048_));
 sky130_fd_sc_hd__or4_2 _0955_ (.A(\Signal_Generator_2_270phase_inst.count[3] ),
    .B(\Signal_Generator_2_270phase_inst.count[2] ),
    .C(\Signal_Generator_2_270phase_inst.count[1] ),
    .D(\Signal_Generator_2_270phase_inst.count[0] ),
    .X(_0422_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(\Signal_Generator_2_270phase_inst.direction ),
    .Y(_0423_));
 sky130_fd_sc_hd__o31a_2 _0957_ (.A1(\Signal_Generator_2_270phase_inst.count[5] ),
    .A2(\Signal_Generator_2_270phase_inst.count[4] ),
    .A3(_0422_),
    .B1(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__and2_1 _0958_ (.A(\Signal_Generator_2_270phase_inst.count[1] ),
    .B(\Signal_Generator_2_270phase_inst.count[0] ),
    .X(_0425_));
 sky130_fd_sc_hd__and3_1 _0959_ (.A(\Signal_Generator_2_270phase_inst.count[3] ),
    .B(\Signal_Generator_2_270phase_inst.count[2] ),
    .C(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__and3_1 _0960_ (.A(\Signal_Generator_2_270phase_inst.count[5] ),
    .B(\Signal_Generator_2_270phase_inst.count[4] ),
    .C(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nor2_1 _0961_ (.A(_0424_),
    .B(_0427_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(net49),
    .Y(_0050_));
 sky130_fd_sc_hd__nor2_1 _0963_ (.A(\Signal_Generator_2_270phase_inst.count[1] ),
    .B(\Signal_Generator_2_270phase_inst.count[0] ),
    .Y(_0428_));
 sky130_fd_sc_hd__or2_1 _0964_ (.A(_0428_),
    .B(_0425_),
    .X(_0429_));
 sky130_fd_sc_hd__a21oi_1 _0965_ (.A1(_0424_),
    .A2(_0429_),
    .B1(\Signal_Generator_2_270phase_inst.direction ),
    .Y(_0430_));
 sky130_fd_sc_hd__a21oi_1 _0966_ (.A1(_0056_),
    .A2(_0429_),
    .B1(_0430_),
    .Y(_0051_));
 sky130_fd_sc_hd__xor2_1 _0967_ (.A(\Signal_Generator_2_270phase_inst.count[2] ),
    .B(_0428_),
    .X(_0431_));
 sky130_fd_sc_hd__xor2_1 _0968_ (.A(\Signal_Generator_2_270phase_inst.count[2] ),
    .B(_0425_),
    .X(_0432_));
 sky130_fd_sc_hd__or2_1 _0969_ (.A(_0427_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _0970_ (.A1(_0424_),
    .A2(_0431_),
    .B1(_0433_),
    .B2(\Signal_Generator_2_270phase_inst.direction ),
    .X(_0052_));
 sky130_fd_sc_hd__o31ai_1 _0971_ (.A1(\Signal_Generator_2_270phase_inst.count[2] ),
    .A2(\Signal_Generator_2_270phase_inst.count[1] ),
    .A3(\Signal_Generator_2_270phase_inst.count[0] ),
    .B1(\Signal_Generator_2_270phase_inst.count[3] ),
    .Y(_0434_));
 sky130_fd_sc_hd__nand2_1 _0972_ (.A(_0422_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_2 _0973_ (.A(_0426_),
    .Y(_0436_));
 sky130_fd_sc_hd__a31o_1 _0974_ (.A1(\Signal_Generator_2_270phase_inst.count[2] ),
    .A2(\Signal_Generator_2_270phase_inst.count[1] ),
    .A3(\Signal_Generator_2_270phase_inst.count[0] ),
    .B1(\Signal_Generator_2_270phase_inst.count[3] ),
    .X(_0437_));
 sky130_fd_sc_hd__a21o_1 _0975_ (.A1(_0436_),
    .A2(_0437_),
    .B1(_0427_),
    .X(_0438_));
 sky130_fd_sc_hd__a22o_1 _0976_ (.A1(_0424_),
    .A2(_0435_),
    .B1(_0438_),
    .B2(\Signal_Generator_2_270phase_inst.direction ),
    .X(_0053_));
 sky130_fd_sc_hd__or3b_1 _0977_ (.A(_0436_),
    .B(\Signal_Generator_2_270phase_inst.count[5] ),
    .C_N(\Signal_Generator_2_270phase_inst.count[4] ),
    .X(_0439_));
 sky130_fd_sc_hd__or2_1 _0978_ (.A(\Signal_Generator_2_270phase_inst.count[4] ),
    .B(_0426_),
    .X(_0440_));
 sky130_fd_sc_hd__xnor2_1 _0979_ (.A(\Signal_Generator_2_270phase_inst.count[4] ),
    .B(_0422_),
    .Y(_0441_));
 sky130_fd_sc_hd__a32o_1 _0980_ (.A1(\Signal_Generator_2_270phase_inst.direction ),
    .A2(_0439_),
    .A3(_0440_),
    .B1(_0424_),
    .B2(_0441_),
    .X(_0054_));
 sky130_fd_sc_hd__o31a_1 _0981_ (.A1(\Signal_Generator_2_270phase_inst.count[4] ),
    .A2(\Signal_Generator_2_270phase_inst.direction ),
    .A3(_0422_),
    .B1(\Signal_Generator_2_270phase_inst.count[5] ),
    .X(_0442_));
 sky130_fd_sc_hd__a31o_1 _0982_ (.A1(\Signal_Generator_2_270phase_inst.count[4] ),
    .A2(\Signal_Generator_2_270phase_inst.direction ),
    .A3(_0426_),
    .B1(_0442_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_2 _0983_ (.A0(CLK_PLL),
    .A1(CLK_EXT),
    .S(\Shift_Register_Inst.data_out[14] ),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_2 _0984_ (.A(_0443_),
    .X(\Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__and2_1 _0985_ (.A(\Shift_Register_Inst.data_out[16] ),
    .B(net8),
    .X(_0444_));
 sky130_fd_sc_hd__buf_1 _0986_ (.A(_0444_),
    .X(net19));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(net41),
    .Y(_0445_));
 sky130_fd_sc_hd__or2_1 _0988_ (.A(_0445_),
    .B(net7),
    .X(_0446_));
 sky130_fd_sc_hd__buf_1 _0989_ (.A(_0446_),
    .X(net24));
 sky130_fd_sc_hd__and3_1 _0990_ (.A(_0445_),
    .B(\Shift_Register_Inst.data_out[17] ),
    .C(NMOS1_PS2_prev),
    .X(_0447_));
 sky130_fd_sc_hd__buf_1 _0991_ (.A(_0447_),
    .X(net16));
 sky130_fd_sc_hd__or2b_1 _0992_ (.A(\Shift_Register_Inst.data_out[16] ),
    .B_N(\Shift_Register_Inst.data_out[17] ),
    .X(_0448_));
 sky130_fd_sc_hd__or2_1 _0993_ (.A(PMOS2_PS2_prev),
    .B(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__buf_1 _0994_ (.A(_0449_),
    .X(net23));
 sky130_fd_sc_hd__and3_1 _0995_ (.A(_0445_),
    .B(\Shift_Register_Inst.data_out[17] ),
    .C(NMOS2_PS2_prev),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _0996_ (.A(_0450_),
    .X(net18));
 sky130_fd_sc_hd__or2_1 _0997_ (.A(PMOS1_PS2_prev),
    .B(_0448_),
    .X(_0451_));
 sky130_fd_sc_hd__buf_1 _0998_ (.A(_0451_),
    .X(net21));
 sky130_fd_sc_hd__and3_1 _0999_ (.A(_0445_),
    .B(\Shift_Register_Inst.data_out[17] ),
    .C(NMOS1_PS1_prev),
    .X(_0452_));
 sky130_fd_sc_hd__buf_1 _1000_ (.A(_0452_),
    .X(net15));
 sky130_fd_sc_hd__or2_1 _1001_ (.A(PMOS2_PS1_prev),
    .B(_0448_),
    .X(_0453_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1002_ (.A(_0453_),
    .X(net22));
 sky130_fd_sc_hd__and3_1 _1003_ (.A(_0445_),
    .B(\Shift_Register_Inst.data_out[17] ),
    .C(NMOS2_PS1_prev),
    .X(_0454_));
 sky130_fd_sc_hd__buf_1 _1004_ (.A(_0454_),
    .X(net17));
 sky130_fd_sc_hd__or2_1 _1005_ (.A(PMOS1_PS1_prev),
    .B(_0448_),
    .X(_0455_));
 sky130_fd_sc_hd__buf_1 _1006_ (.A(_0455_),
    .X(net20));
 sky130_fd_sc_hd__and2b_1 _1007_ (.A_N(\Shift_Register_Inst.data_out[10] ),
    .B(\Shift_Register_Inst.data_out[9] ),
    .X(_0456_));
 sky130_fd_sc_hd__and2_1 _1008_ (.A(net19),
    .B(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__nor2_1 _1009_ (.A(\Shift_Register_Inst.data_out[9] ),
    .B(\Shift_Register_Inst.data_out[10] ),
    .Y(_0458_));
 sky130_fd_sc_hd__and2b_1 _1010_ (.A_N(\Shift_Register_Inst.data_out[9] ),
    .B(\Shift_Register_Inst.data_out[10] ),
    .X(_0459_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(\Shift_Register_Inst.data_out[12] ),
    .Y(_0460_));
 sky130_fd_sc_hd__a221o_2 _1012_ (.A1(net24),
    .A2(_0458_),
    .B1(_0459_),
    .B2(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ),
    .C1(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__a211o_1 _1013_ (.A1(net20),
    .A2(_0458_),
    .B1(\Shift_Register_Inst.data_out[11] ),
    .C1(\Shift_Register_Inst.data_out[12] ),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _1014_ (.A1(net17),
    .A2(_0456_),
    .B1(_0459_),
    .B2(net22),
    .X(_0463_));
 sky130_fd_sc_hd__a31o_1 _1015_ (.A1(\Shift_Register_Inst.data_out[9] ),
    .A2(\Shift_Register_Inst.data_out[10] ),
    .A3(net15),
    .B1(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__or2_1 _1016_ (.A(_0462_),
    .B(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__and2_1 _1017_ (.A(_0445_),
    .B(\Shift_Register_Inst.data_out[17] ),
    .X(_0466_));
 sky130_fd_sc_hd__and3_1 _1018_ (.A(NMOS2_PS2_prev),
    .B(_0466_),
    .C(_0456_),
    .X(_0467_));
 sky130_fd_sc_hd__and2_1 _1019_ (.A(net21),
    .B(_0458_),
    .X(_0468_));
 sky130_fd_sc_hd__a31o_1 _1020_ (.A1(\Shift_Register_Inst.data_out[9] ),
    .A2(\Shift_Register_Inst.data_out[10] ),
    .A3(net16),
    .B1(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a211oi_1 _1021_ (.A1(net23),
    .A2(_0459_),
    .B1(_0467_),
    .C1(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__o21ai_1 _1022_ (.A1(\Shift_Register_Inst.data_out[12] ),
    .A2(_0470_),
    .B1(\Shift_Register_Inst.data_out[11] ),
    .Y(_0471_));
 sky130_fd_sc_hd__o211a_4 _1023_ (.A1(_0457_),
    .A2(_0461_),
    .B1(_0465_),
    .C1(_0471_),
    .X(net25));
 sky130_fd_sc_hd__nand2_1 _1024_ (.A(_0262_),
    .B(net6),
    .Y(_0472_));
 sky130_fd_sc_hd__o211ai_1 _1025_ (.A1(_0262_),
    .A2(\Dead_Time_Generator_inst_1.go ),
    .B1(_0472_),
    .C1(net31),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_1 _1026_ (.A(_0262_),
    .B(net4),
    .Y(_0473_));
 sky130_fd_sc_hd__o211ai_1 _1027_ (.A1(_0262_),
    .A2(\Dead_Time_Generator_inst_3.go ),
    .B1(_0473_),
    .C1(net31),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(net31),
    .Y(_0474_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(\Dead_Time_Generator_inst_2.go ),
    .A1(net3),
    .S(_0262_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _1030_ (.A(_0474_),
    .B(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0476_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(\Dead_Time_Generator_inst_4.go ),
    .A1(net5),
    .S(_0262_),
    .X(_0477_));
 sky130_fd_sc_hd__and2_1 _1033_ (.A(_0474_),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(_0478_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _1035_ (.A(net31),
    .B(_0475_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(_0479_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1037_ (.A(net31),
    .B(_0477_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(_0480_),
    .X(_0000_));
 sky130_fd_sc_hd__o211ai_1 _1039_ (.A1(_0262_),
    .A2(net36),
    .B1(_0472_),
    .C1(_0474_),
    .Y(_0005_));
 sky130_fd_sc_hd__o211ai_1 _1040_ (.A1(_0262_),
    .A2(net35),
    .B1(_0473_),
    .C1(_0474_),
    .Y(_0007_));
 sky130_fd_sc_hd__buf_2 _1041_ (.A(net2),
    .X(_0481_));
 sky130_fd_sc_hd__buf_4 _1042_ (.A(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_4 _1043_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__inv_2 _1044_ (.A(_0483_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(_0483_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(_0483_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(_0483_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(_0483_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(_0483_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(_0483_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(_0483_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(_0483_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(_0483_),
    .Y(_0073_));
 sky130_fd_sc_hd__buf_4 _1054_ (.A(_0482_),
    .X(_0484_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(_0484_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(_0484_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(_0484_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0484_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(_0484_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(_0484_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(_0484_),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0484_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0484_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(_0484_),
    .Y(_0083_));
 sky130_fd_sc_hd__buf_4 _1065_ (.A(_0482_),
    .X(_0485_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(_0485_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(_0485_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(_0485_),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(_0485_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0485_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(_0485_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(_0485_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0485_),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(_0485_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(_0485_),
    .Y(_0093_));
 sky130_fd_sc_hd__or2b_1 _1076_ (.A(net37),
    .B_N(\Dead_Time_Generator_inst_4.count_dt[4] ),
    .X(_0486_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(\Dead_Time_Generator_inst_4.count_dt[3] ),
    .Y(_0487_));
 sky130_fd_sc_hd__inv_2 _1078_ (.A(\Dead_Time_Generator_inst_4.count_dt[0] ),
    .Y(_0488_));
 sky130_fd_sc_hd__or2b_1 _1079_ (.A(\Dead_Time_Generator_inst_1.dt[1] ),
    .B_N(\Dead_Time_Generator_inst_4.count_dt[1] ),
    .X(_0489_));
 sky130_fd_sc_hd__and2b_1 _1080_ (.A_N(\Dead_Time_Generator_inst_4.count_dt[2] ),
    .B(\Dead_Time_Generator_inst_1.dt[2] ),
    .X(_0490_));
 sky130_fd_sc_hd__and2b_1 _1081_ (.A_N(\Dead_Time_Generator_inst_4.count_dt[1] ),
    .B(\Dead_Time_Generator_inst_1.dt[1] ),
    .X(_0491_));
 sky130_fd_sc_hd__a311o_1 _1082_ (.A1(_0488_),
    .A2(\Dead_Time_Generator_inst_1.dt[0] ),
    .A3(_0489_),
    .B1(_0490_),
    .C1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(\Dead_Time_Generator_inst_4.count_dt[2] ),
    .Y(_0493_));
 sky130_fd_sc_hd__o22a_1 _1084_ (.A1(_0493_),
    .A2(\Dead_Time_Generator_inst_1.dt[2] ),
    .B1(net45),
    .B2(_0487_),
    .X(_0494_));
 sky130_fd_sc_hd__and2b_1 _1085_ (.A_N(\Dead_Time_Generator_inst_4.count_dt[4] ),
    .B(net37),
    .X(_0495_));
 sky130_fd_sc_hd__a221o_1 _1086_ (.A1(_0487_),
    .A2(net39),
    .B1(_0492_),
    .B2(net46),
    .C1(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__nand2_1 _1087_ (.A(_0486_),
    .B(net47),
    .Y(_0497_));
 sky130_fd_sc_hd__or2_1 _1088_ (.A(_0248_),
    .B(_0250_),
    .X(_0498_));
 sky130_fd_sc_hd__and2b_1 _1089_ (.A_N(\Shift_Register_Inst.data_out[7] ),
    .B(\Shift_Register_Inst.data_out[8] ),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_1 _1090_ (.A(\Shift_Register_Inst.data_out[7] ),
    .B(_0250_),
    .Y(_0500_));
 sky130_fd_sc_hd__and3_1 _1091_ (.A(\Shift_Register_Inst.data_out[7] ),
    .B(\Shift_Register_Inst.data_out[8] ),
    .C(\Signal_Generator_2_270phase_inst.count[4] ),
    .X(_0501_));
 sky130_fd_sc_hd__and3b_1 _1092_ (.A_N(\Shift_Register_Inst.data_out[8] ),
    .B(\Signal_Generator_2_90phase_inst.count[4] ),
    .C(_0248_),
    .X(_0502_));
 sky130_fd_sc_hd__a2111o_1 _1093_ (.A1(\Signal_Generator_2_180phase_inst.count[4] ),
    .A2(_0499_),
    .B1(_0500_),
    .C1(_0501_),
    .D1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o21ai_1 _1094_ (.A1(\Signal_Generator_2_0phase_inst.count[4] ),
    .A2(_0498_),
    .B1(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(net14),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _1096_ (.A(\Shift_Register_Inst.data_out[8] ),
    .Y(_0506_));
 sky130_fd_sc_hd__and3_1 _1097_ (.A(_0248_),
    .B(_0506_),
    .C(\Signal_Generator_2_90phase_inst.count[5] ),
    .X(_0507_));
 sky130_fd_sc_hd__and3_1 _1098_ (.A(_0248_),
    .B(_0250_),
    .C(\Signal_Generator_2_270phase_inst.count[5] ),
    .X(_0508_));
 sky130_fd_sc_hd__a21o_1 _1099_ (.A1(\Signal_Generator_2_180phase_inst.count[5] ),
    .A2(_0499_),
    .B1(_0500_),
    .X(_0509_));
 sky130_fd_sc_hd__o32a_1 _1100_ (.A1(_0507_),
    .A2(_0508_),
    .A3(_0509_),
    .B1(_0498_),
    .B2(\Signal_Generator_2_0phase_inst.count[5] ),
    .X(_0510_));
 sky130_fd_sc_hd__a2bb2o_1 _1101_ (.A1_N(_0504_),
    .A2_N(net13),
    .B1(_0505_),
    .B2(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__or2_1 _1102_ (.A(_0505_),
    .B(_0510_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_1 _1103_ (.A(net13),
    .B(_0504_),
    .Y(_0513_));
 sky130_fd_sc_hd__and3b_1 _1104_ (.A_N(_0511_),
    .B(_0512_),
    .C(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__inv_2 _1105_ (.A(net12),
    .Y(_0515_));
 sky130_fd_sc_hd__and3b_1 _1106_ (.A_N(\Shift_Register_Inst.data_out[8] ),
    .B(\Signal_Generator_2_90phase_inst.count[3] ),
    .C(\Shift_Register_Inst.data_out[7] ),
    .X(_0516_));
 sky130_fd_sc_hd__and3_1 _1107_ (.A(\Shift_Register_Inst.data_out[7] ),
    .B(\Shift_Register_Inst.data_out[8] ),
    .C(\Signal_Generator_2_270phase_inst.count[3] ),
    .X(_0517_));
 sky130_fd_sc_hd__and3b_1 _1108_ (.A_N(\Shift_Register_Inst.data_out[7] ),
    .B(\Shift_Register_Inst.data_out[8] ),
    .C(\Signal_Generator_2_180phase_inst.count[3] ),
    .X(_0518_));
 sky130_fd_sc_hd__or4_1 _1109_ (.A(_0500_),
    .B(_0516_),
    .C(_0517_),
    .D(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _1110_ (.A(\Signal_Generator_2_0phase_inst.count[3] ),
    .B(_0498_),
    .X(_0520_));
 sky130_fd_sc_hd__and3_1 _1111_ (.A(_0515_),
    .B(_0519_),
    .C(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__inv_2 _1112_ (.A(net11),
    .Y(_0522_));
 sky130_fd_sc_hd__and3b_1 _1113_ (.A_N(\Shift_Register_Inst.data_out[7] ),
    .B(_0250_),
    .C(\Signal_Generator_2_180phase_inst.count[2] ),
    .X(_0523_));
 sky130_fd_sc_hd__and3_1 _1114_ (.A(_0248_),
    .B(_0250_),
    .C(\Signal_Generator_2_270phase_inst.count[2] ),
    .X(_0524_));
 sky130_fd_sc_hd__a2111o_1 _1115_ (.A1(_0506_),
    .A2(\Signal_Generator_2_90phase_inst.count[2] ),
    .B1(_0500_),
    .C1(_0523_),
    .D1(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_1 _1116_ (.A(\Signal_Generator_2_0phase_inst.count[2] ),
    .B(_0498_),
    .X(_0526_));
 sky130_fd_sc_hd__and3_1 _1117_ (.A(_0522_),
    .B(_0525_),
    .C(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__a21o_1 _1118_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0515_),
    .X(_0528_));
 sky130_fd_sc_hd__a21o_1 _1119_ (.A1(_0525_),
    .A2(_0526_),
    .B1(_0522_),
    .X(_0529_));
 sky130_fd_sc_hd__and4bb_1 _1120_ (.A_N(_0521_),
    .B_N(_0527_),
    .C(_0528_),
    .D(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__or2_1 _1121_ (.A(\Signal_Generator_2_0phase_inst.count[1] ),
    .B(_0498_),
    .X(_0531_));
 sky130_fd_sc_hd__and3b_1 _1122_ (.A_N(_0250_),
    .B(\Signal_Generator_2_90phase_inst.count[1] ),
    .C(_0248_),
    .X(_0532_));
 sky130_fd_sc_hd__and3b_1 _1123_ (.A_N(_0248_),
    .B(_0250_),
    .C(\Signal_Generator_2_180phase_inst.count[1] ),
    .X(_0533_));
 sky130_fd_sc_hd__and3_1 _1124_ (.A(_0248_),
    .B(_0250_),
    .C(\Signal_Generator_2_270phase_inst.count[1] ),
    .X(_0534_));
 sky130_fd_sc_hd__or4_1 _1125_ (.A(_0500_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(net10),
    .Y(_0536_));
 sky130_fd_sc_hd__a21o_1 _1127_ (.A1(_0531_),
    .A2(_0535_),
    .B1(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__mux4_1 _1128_ (.A0(\Signal_Generator_2_0phase_inst.count[0] ),
    .A1(\Signal_Generator_2_90phase_inst.count[0] ),
    .A2(\Signal_Generator_2_180phase_inst.count[0] ),
    .A3(\Signal_Generator_2_270phase_inst.count[0] ),
    .S0(_0248_),
    .S1(_0250_),
    .X(_0538_));
 sky130_fd_sc_hd__or2b_1 _1129_ (.A(_0538_),
    .B_N(net9),
    .X(_0539_));
 sky130_fd_sc_hd__and3_1 _1130_ (.A(_0536_),
    .B(_0531_),
    .C(_0535_),
    .X(_0540_));
 sky130_fd_sc_hd__a21o_1 _1131_ (.A1(_0537_),
    .A2(_0539_),
    .B1(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__o21a_1 _1132_ (.A1(_0521_),
    .A2(_0527_),
    .B1(_0528_),
    .X(_0542_));
 sky130_fd_sc_hd__a21o_1 _1133_ (.A1(_0530_),
    .A2(_0541_),
    .B1(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _1134_ (.A1(_0511_),
    .A2(_0512_),
    .B1(_0514_),
    .B2(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__buf_2 _1135_ (.A(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__and2b_1 _1136_ (.A_N(net9),
    .B(_0538_),
    .X(_0546_));
 sky130_fd_sc_hd__nand3b_1 _1137_ (.A_N(_0540_),
    .B(_0537_),
    .C(_0539_),
    .Y(_0547_));
 sky130_fd_sc_hd__or4bb_2 _1138_ (.A(_0546_),
    .B(_0547_),
    .C_N(_0530_),
    .D_N(_0514_),
    .X(_0548_));
 sky130_fd_sc_hd__buf_2 _1139_ (.A(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__and3_1 _1140_ (.A(_0497_),
    .B(_0545_),
    .C(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_1 _1141_ (.A(_0550_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_4 _1142_ (.A(_0481_),
    .X(_0551_));
 sky130_fd_sc_hd__inv_2 _1143_ (.A(_0551_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1144_ (.A(_0551_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1145_ (.A(_0551_),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1146_ (.A(_0551_),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1147_ (.A(_0551_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1148_ (.A(_0551_),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _1149_ (.A(_0551_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1150_ (.A(_0551_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1151_ (.A(_0551_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1152_ (.A(_0551_),
    .Y(_0103_));
 sky130_fd_sc_hd__buf_4 _1153_ (.A(_0481_),
    .X(_0552_));
 sky130_fd_sc_hd__inv_2 _1154_ (.A(_0552_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1155_ (.A(_0552_),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1156_ (.A(_0552_),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1157_ (.A(_0552_),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1158_ (.A(_0552_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1159_ (.A(_0552_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _1160_ (.A(_0552_),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1161_ (.A(_0552_),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _1162_ (.A(_0552_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1163_ (.A(_0552_),
    .Y(_0113_));
 sky130_fd_sc_hd__buf_4 _1164_ (.A(_0481_),
    .X(_0553_));
 sky130_fd_sc_hd__inv_2 _1165_ (.A(_0553_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1166_ (.A(_0553_),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1167_ (.A(_0553_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1168_ (.A(_0553_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(_0553_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1170_ (.A(_0553_),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1171_ (.A(_0553_),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1172_ (.A(_0553_),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1173_ (.A(_0553_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1174_ (.A(_0553_),
    .Y(_0123_));
 sky130_fd_sc_hd__buf_4 _1175_ (.A(_0481_),
    .X(_0554_));
 sky130_fd_sc_hd__inv_2 _1176_ (.A(_0554_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1177_ (.A(_0554_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1178_ (.A(_0554_),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1179_ (.A(_0554_),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1180_ (.A(_0554_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1181_ (.A(_0554_),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1182_ (.A(_0554_),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1183_ (.A(_0554_),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1184_ (.A(_0554_),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1185_ (.A(_0554_),
    .Y(_0133_));
 sky130_fd_sc_hd__buf_4 _1186_ (.A(_0481_),
    .X(_0555_));
 sky130_fd_sc_hd__inv_2 _1187_ (.A(_0555_),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1188_ (.A(_0555_),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1189_ (.A(_0555_),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1190_ (.A(_0555_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1191_ (.A(_0555_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1192_ (.A(_0555_),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(_0555_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1194_ (.A(_0555_),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1195_ (.A(_0555_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1196_ (.A(_0555_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1197_ (.A(_0482_),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1198_ (.A(_0482_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1199_ (.A(_0482_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1200_ (.A(_0482_),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(_0482_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1202_ (.A(_0482_),
    .Y(_0149_));
 sky130_fd_sc_hd__nand2_1 _1203_ (.A(_0445_),
    .B(net8),
    .Y(_0556_));
 sky130_fd_sc_hd__clkbuf_2 _1204_ (.A(\Shift_Register_Inst.data_out[6] ),
    .X(_0557_));
 sky130_fd_sc_hd__or2_1 _1205_ (.A(_0242_),
    .B(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__and3b_1 _1206_ (.A_N(_0242_),
    .B(_0245_),
    .C(\Signal_Generator_1_180phase_inst.count[5] ),
    .X(_0559_));
 sky130_fd_sc_hd__a31o_1 _1207_ (.A1(_0242_),
    .A2(_0245_),
    .A3(\Signal_Generator_1_270phase_inst.count[5] ),
    .B1(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _1208_ (.A1(_0242_),
    .A2(_0312_),
    .B1(_0245_),
    .Y(_0561_));
 sky130_fd_sc_hd__o22a_1 _1209_ (.A1(\Signal_Generator_1_0phase_inst.count[5] ),
    .A2(_0558_),
    .B1(_0560_),
    .B2(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__nor2_1 _1210_ (.A(_0556_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_2 _1211_ (.A(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _1212_ (.A(_0445_),
    .B(net7),
    .Y(_0565_));
 sky130_fd_sc_hd__and3_1 _1213_ (.A(_0242_),
    .B(_0245_),
    .C(\Signal_Generator_1_270phase_inst.count[4] ),
    .X(_0566_));
 sky130_fd_sc_hd__inv_2 _1214_ (.A(_0245_),
    .Y(_0567_));
 sky130_fd_sc_hd__nor2_2 _1215_ (.A(_0241_),
    .B(\Shift_Register_Inst.data_out[6] ),
    .Y(_0568_));
 sky130_fd_sc_hd__and3b_1 _1216_ (.A_N(_0242_),
    .B(_0245_),
    .C(\Signal_Generator_1_180phase_inst.count[4] ),
    .X(_0569_));
 sky130_fd_sc_hd__a211o_1 _1217_ (.A1(_0567_),
    .A2(\Signal_Generator_1_90phase_inst.count[4] ),
    .B1(_0568_),
    .C1(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__o22a_1 _1218_ (.A1(\Signal_Generator_1_0phase_inst.count[4] ),
    .A2(_0558_),
    .B1(_0566_),
    .B2(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__a22o_1 _1219_ (.A1(_0556_),
    .A2(_0562_),
    .B1(_0565_),
    .B2(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__or2_1 _1220_ (.A(\Signal_Generator_1_0phase_inst.count[1] ),
    .B(_0558_),
    .X(_0573_));
 sky130_fd_sc_hd__and3b_1 _1221_ (.A_N(\Shift_Register_Inst.data_out[5] ),
    .B(\Shift_Register_Inst.data_out[6] ),
    .C(\Signal_Generator_1_180phase_inst.count[1] ),
    .X(_0574_));
 sky130_fd_sc_hd__and3b_1 _1222_ (.A_N(\Shift_Register_Inst.data_out[6] ),
    .B(\Signal_Generator_1_90phase_inst.count[1] ),
    .C(_0241_),
    .X(_0575_));
 sky130_fd_sc_hd__and3_1 _1223_ (.A(_0241_),
    .B(_0557_),
    .C(\Signal_Generator_1_270phase_inst.count[1] ),
    .X(_0576_));
 sky130_fd_sc_hd__or4_1 _1224_ (.A(_0568_),
    .B(_0574_),
    .C(_0575_),
    .D(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__inv_2 _1225_ (.A(net4),
    .Y(_0578_));
 sky130_fd_sc_hd__a211o_1 _1226_ (.A1(_0573_),
    .A2(_0577_),
    .B1(net33),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__and3b_1 _1227_ (.A_N(_0241_),
    .B(_0557_),
    .C(\Signal_Generator_1_180phase_inst.count[0] ),
    .X(_0580_));
 sky130_fd_sc_hd__and3b_1 _1228_ (.A_N(_0557_),
    .B(\Signal_Generator_1_90phase_inst.count[0] ),
    .C(_0241_),
    .X(_0581_));
 sky130_fd_sc_hd__and3_1 _1229_ (.A(_0242_),
    .B(_0245_),
    .C(\Signal_Generator_1_270phase_inst.count[0] ),
    .X(_0582_));
 sky130_fd_sc_hd__or4_1 _1230_ (.A(_0568_),
    .B(_0580_),
    .C(_0581_),
    .D(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _1231_ (.A(_0008_),
    .B(_0568_),
    .Y(_0584_));
 sky130_fd_sc_hd__or2b_1 _1232_ (.A(net33),
    .B_N(net3),
    .X(_0585_));
 sky130_fd_sc_hd__a21o_1 _1233_ (.A1(_0583_),
    .A2(_0584_),
    .B1(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__o211a_1 _1234_ (.A1(_0262_),
    .A2(_0578_),
    .B1(_0573_),
    .C1(_0577_),
    .X(_0587_));
 sky130_fd_sc_hd__a21o_1 _1235_ (.A1(_0579_),
    .A2(_0586_),
    .B1(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__or2b_1 _1236_ (.A(net33),
    .B_N(net6),
    .X(_0589_));
 sky130_fd_sc_hd__and3_1 _1237_ (.A(_0241_),
    .B(_0557_),
    .C(\Signal_Generator_1_270phase_inst.count[3] ),
    .X(_0590_));
 sky130_fd_sc_hd__and3b_1 _1238_ (.A_N(_0241_),
    .B(_0557_),
    .C(\Signal_Generator_1_180phase_inst.count[3] ),
    .X(_0591_));
 sky130_fd_sc_hd__and2b_1 _1239_ (.A_N(_0557_),
    .B(\Signal_Generator_1_90phase_inst.count[3] ),
    .X(_0592_));
 sky130_fd_sc_hd__or3_1 _1240_ (.A(_0242_),
    .B(_0245_),
    .C(\Signal_Generator_1_0phase_inst.count[3] ),
    .X(_0593_));
 sky130_fd_sc_hd__o41a_1 _1241_ (.A1(_0568_),
    .A2(_0590_),
    .A3(_0591_),
    .A4(_0592_),
    .B1(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__or2b_1 _1242_ (.A(net33),
    .B_N(net5),
    .X(_0595_));
 sky130_fd_sc_hd__and3_1 _1243_ (.A(_0241_),
    .B(_0557_),
    .C(\Signal_Generator_1_270phase_inst.count[2] ),
    .X(_0596_));
 sky130_fd_sc_hd__and3b_1 _1244_ (.A_N(_0241_),
    .B(_0557_),
    .C(\Signal_Generator_1_180phase_inst.count[2] ),
    .X(_0597_));
 sky130_fd_sc_hd__and2b_1 _1245_ (.A_N(_0557_),
    .B(\Signal_Generator_1_90phase_inst.count[2] ),
    .X(_0598_));
 sky130_fd_sc_hd__or3_1 _1246_ (.A(_0242_),
    .B(_0245_),
    .C(\Signal_Generator_1_0phase_inst.count[2] ),
    .X(_0599_));
 sky130_fd_sc_hd__o41a_1 _1247_ (.A1(_0568_),
    .A2(_0596_),
    .A3(_0597_),
    .A4(_0598_),
    .B1(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__o22a_1 _1248_ (.A1(_0589_),
    .A2(_0594_),
    .B1(_0595_),
    .B2(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__a22o_1 _1249_ (.A1(_0589_),
    .A2(_0594_),
    .B1(_0595_),
    .B2(_0600_),
    .X(_0602_));
 sky130_fd_sc_hd__o21a_1 _1250_ (.A1(_0589_),
    .A2(_0594_),
    .B1(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_1 _1251_ (.A1(_0588_),
    .A2(_0601_),
    .B1(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _1252_ (.A(_0565_),
    .B(_0571_),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _1253_ (.A(_0563_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__a22o_1 _1254_ (.A1(_0564_),
    .A2(_0572_),
    .B1(_0604_),
    .B2(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__and3_1 _1255_ (.A(_0583_),
    .B(_0584_),
    .C(_0585_),
    .X(_0608_));
 sky130_fd_sc_hd__or4bb_1 _1256_ (.A(_0602_),
    .B(_0587_),
    .C_N(_0579_),
    .D_N(_0586_),
    .X(_0609_));
 sky130_fd_sc_hd__or4_1 _1257_ (.A(_0563_),
    .B(_0572_),
    .C(_0605_),
    .D(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__or3b_1 _1258_ (.A(_0608_),
    .B(_0610_),
    .C_N(_0601_),
    .X(_0611_));
 sky130_fd_sc_hd__or2b_1 _1259_ (.A(net37),
    .B_N(\Dead_Time_Generator_inst_1.count_dt[4] ),
    .X(_0612_));
 sky130_fd_sc_hd__inv_2 _1260_ (.A(net54),
    .Y(_0613_));
 sky130_fd_sc_hd__inv_2 _1261_ (.A(net70),
    .Y(_0614_));
 sky130_fd_sc_hd__or2b_1 _1262_ (.A(\Dead_Time_Generator_inst_1.dt[1] ),
    .B_N(\Dead_Time_Generator_inst_1.count_dt[1] ),
    .X(_0615_));
 sky130_fd_sc_hd__and2b_1 _1263_ (.A_N(\Dead_Time_Generator_inst_1.count_dt[0] ),
    .B(\Dead_Time_Generator_inst_1.dt[0] ),
    .X(_0616_));
 sky130_fd_sc_hd__and2b_1 _1264_ (.A_N(\Dead_Time_Generator_inst_1.count_dt[1] ),
    .B(\Dead_Time_Generator_inst_1.dt[1] ),
    .X(_0617_));
 sky130_fd_sc_hd__a221o_1 _1265_ (.A1(_0614_),
    .A2(\Dead_Time_Generator_inst_1.dt[2] ),
    .B1(_0615_),
    .B2(_0616_),
    .C1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__o22a_1 _1266_ (.A1(_0614_),
    .A2(\Dead_Time_Generator_inst_1.dt[2] ),
    .B1(net39),
    .B2(_0613_),
    .X(_0619_));
 sky130_fd_sc_hd__and2b_1 _1267_ (.A_N(\Dead_Time_Generator_inst_1.count_dt[4] ),
    .B(net37),
    .X(_0620_));
 sky130_fd_sc_hd__a221o_1 _1268_ (.A1(_0613_),
    .A2(net39),
    .B1(_0618_),
    .B2(_0619_),
    .C1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__and3_1 _1269_ (.A(\Dead_Time_Generator_inst_1.count_dt[0] ),
    .B(_0612_),
    .C(net40),
    .X(_0622_));
 sky130_fd_sc_hd__and2_1 _1270_ (.A(_0612_),
    .B(net40),
    .X(_0623_));
 sky130_fd_sc_hd__nor2_1 _1271_ (.A(\Dead_Time_Generator_inst_1.count_dt[0] ),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__a211oi_1 _1272_ (.A1(_0607_),
    .A2(_0611_),
    .B1(_0622_),
    .C1(_0624_),
    .Y(_0174_));
 sky130_fd_sc_hd__buf_2 _1273_ (.A(_0607_),
    .X(_0625_));
 sky130_fd_sc_hd__buf_2 _1274_ (.A(_0611_),
    .X(_0626_));
 sky130_fd_sc_hd__nand2_1 _1275_ (.A(\Dead_Time_Generator_inst_1.count_dt[1] ),
    .B(_0622_),
    .Y(_0627_));
 sky130_fd_sc_hd__or2_1 _1276_ (.A(\Dead_Time_Generator_inst_1.count_dt[1] ),
    .B(_0622_),
    .X(_0628_));
 sky130_fd_sc_hd__nand2_1 _1277_ (.A(_0627_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__a21oi_1 _1278_ (.A1(_0625_),
    .A2(_0626_),
    .B1(_0629_),
    .Y(_0175_));
 sky130_fd_sc_hd__xnor2_1 _1279_ (.A(_0614_),
    .B(_0627_),
    .Y(_0630_));
 sky130_fd_sc_hd__a21oi_1 _1280_ (.A1(_0625_),
    .A2(_0626_),
    .B1(_0630_),
    .Y(_0176_));
 sky130_fd_sc_hd__and4_1 _1281_ (.A(\Dead_Time_Generator_inst_1.count_dt[3] ),
    .B(\Dead_Time_Generator_inst_1.count_dt[2] ),
    .C(\Dead_Time_Generator_inst_1.count_dt[1] ),
    .D(_0622_),
    .X(_0631_));
 sky130_fd_sc_hd__o21a_1 _1282_ (.A1(_0614_),
    .A2(_0627_),
    .B1(_0613_),
    .X(_0632_));
 sky130_fd_sc_hd__a211oi_1 _1283_ (.A1(_0607_),
    .A2(_0611_),
    .B1(_0631_),
    .C1(_0632_),
    .Y(_0177_));
 sky130_fd_sc_hd__o2bb2a_1 _1284_ (.A1_N(_0625_),
    .A2_N(_0626_),
    .B1(_0631_),
    .B2(net50),
    .X(_0178_));
 sky130_fd_sc_hd__inv_2 _1285_ (.A(_0482_),
    .Y(_0150_));
 sky130_fd_sc_hd__or2b_1 _1286_ (.A(net37),
    .B_N(\Dead_Time_Generator_inst_2.count_dt[4] ),
    .X(_0633_));
 sky130_fd_sc_hd__inv_2 _1287_ (.A(\Dead_Time_Generator_inst_2.count_dt[3] ),
    .Y(_0634_));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(\Dead_Time_Generator_inst_2.count_dt[0] ),
    .Y(_0635_));
 sky130_fd_sc_hd__or2b_1 _1289_ (.A(\Dead_Time_Generator_inst_1.dt[1] ),
    .B_N(\Dead_Time_Generator_inst_2.count_dt[1] ),
    .X(_0636_));
 sky130_fd_sc_hd__and2b_1 _1290_ (.A_N(\Dead_Time_Generator_inst_2.count_dt[2] ),
    .B(\Dead_Time_Generator_inst_1.dt[2] ),
    .X(_0637_));
 sky130_fd_sc_hd__and2b_1 _1291_ (.A_N(\Dead_Time_Generator_inst_2.count_dt[1] ),
    .B(\Dead_Time_Generator_inst_1.dt[1] ),
    .X(_0638_));
 sky130_fd_sc_hd__a311o_1 _1292_ (.A1(_0635_),
    .A2(\Dead_Time_Generator_inst_1.dt[0] ),
    .A3(_0636_),
    .B1(_0637_),
    .C1(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__inv_2 _1293_ (.A(\Dead_Time_Generator_inst_2.count_dt[2] ),
    .Y(_0640_));
 sky130_fd_sc_hd__o22a_1 _1294_ (.A1(_0640_),
    .A2(\Dead_Time_Generator_inst_1.dt[2] ),
    .B1(net45),
    .B2(_0634_),
    .X(_0641_));
 sky130_fd_sc_hd__and2b_1 _1295_ (.A_N(\Dead_Time_Generator_inst_2.count_dt[4] ),
    .B(net53),
    .X(_0642_));
 sky130_fd_sc_hd__a221o_1 _1296_ (.A1(_0634_),
    .A2(net39),
    .B1(_0639_),
    .B2(_0641_),
    .C1(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _1297_ (.A(\Dead_Time_Generator_inst_2.count_dt[0] ),
    .B(_0633_),
    .C(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0633_),
    .B(_0643_),
    .Y(_0645_));
 sky130_fd_sc_hd__and2_1 _1299_ (.A(_0635_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__nor2_1 _1300_ (.A(_0644_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__and3_1 _1301_ (.A(_0625_),
    .B(_0626_),
    .C(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_1 _1302_ (.A(_0648_),
    .X(_0180_));
 sky130_fd_sc_hd__xor2_1 _1303_ (.A(\Dead_Time_Generator_inst_2.count_dt[1] ),
    .B(_0644_),
    .X(_0649_));
 sky130_fd_sc_hd__and3_1 _1304_ (.A(_0625_),
    .B(_0626_),
    .C(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_1 _1305_ (.A(_0650_),
    .X(_0181_));
 sky130_fd_sc_hd__and3_1 _1306_ (.A(\Dead_Time_Generator_inst_2.count_dt[2] ),
    .B(\Dead_Time_Generator_inst_2.count_dt[1] ),
    .C(_0644_),
    .X(_0651_));
 sky130_fd_sc_hd__a21o_1 _1307_ (.A1(\Dead_Time_Generator_inst_2.count_dt[1] ),
    .A2(_0644_),
    .B1(\Dead_Time_Generator_inst_2.count_dt[2] ),
    .X(_0652_));
 sky130_fd_sc_hd__and2b_1 _1308_ (.A_N(_0651_),
    .B(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__and3_1 _1309_ (.A(_0625_),
    .B(_0626_),
    .C(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__clkbuf_1 _1310_ (.A(_0654_),
    .X(_0182_));
 sky130_fd_sc_hd__xnor2_1 _1311_ (.A(_0634_),
    .B(_0651_),
    .Y(_0655_));
 sky130_fd_sc_hd__and3_1 _1312_ (.A(_0625_),
    .B(_0626_),
    .C(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_1 _1313_ (.A(_0656_),
    .X(_0183_));
 sky130_fd_sc_hd__a21o_1 _1314_ (.A1(\Dead_Time_Generator_inst_2.count_dt[3] ),
    .A2(_0651_),
    .B1(\Dead_Time_Generator_inst_2.count_dt[4] ),
    .X(_0657_));
 sky130_fd_sc_hd__and3_1 _1315_ (.A(_0625_),
    .B(_0626_),
    .C(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_1 _1316_ (.A(_0658_),
    .X(_0184_));
 sky130_fd_sc_hd__a21oi_1 _1317_ (.A1(_0625_),
    .A2(_0626_),
    .B1(_0623_),
    .Y(_0185_));
 sky130_fd_sc_hd__or2b_1 _1318_ (.A(net37),
    .B_N(\Dead_Time_Generator_inst_3.count_dt[4] ),
    .X(_0659_));
 sky130_fd_sc_hd__inv_2 _1319_ (.A(net71),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _1320_ (.A(net74),
    .Y(_0661_));
 sky130_fd_sc_hd__or2b_1 _1321_ (.A(\Dead_Time_Generator_inst_1.dt[1] ),
    .B_N(\Dead_Time_Generator_inst_3.count_dt[1] ),
    .X(_0662_));
 sky130_fd_sc_hd__and2b_1 _1322_ (.A_N(\Dead_Time_Generator_inst_3.count_dt[0] ),
    .B(\Dead_Time_Generator_inst_1.dt[0] ),
    .X(_0663_));
 sky130_fd_sc_hd__and2b_1 _1323_ (.A_N(\Dead_Time_Generator_inst_3.count_dt[1] ),
    .B(\Dead_Time_Generator_inst_1.dt[1] ),
    .X(_0664_));
 sky130_fd_sc_hd__a221o_1 _1324_ (.A1(_0661_),
    .A2(\Dead_Time_Generator_inst_1.dt[2] ),
    .B1(_0662_),
    .B2(_0663_),
    .C1(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__o22a_1 _1325_ (.A1(_0661_),
    .A2(\Dead_Time_Generator_inst_1.dt[2] ),
    .B1(net39),
    .B2(_0660_),
    .X(_0666_));
 sky130_fd_sc_hd__and2b_1 _1326_ (.A_N(\Dead_Time_Generator_inst_3.count_dt[4] ),
    .B(net37),
    .X(_0667_));
 sky130_fd_sc_hd__a221o_1 _1327_ (.A1(_0660_),
    .A2(net39),
    .B1(_0665_),
    .B2(_0666_),
    .C1(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__and3_1 _1328_ (.A(\Dead_Time_Generator_inst_3.count_dt[0] ),
    .B(_0659_),
    .C(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__and2_1 _1329_ (.A(_0659_),
    .B(_0668_),
    .X(_0670_));
 sky130_fd_sc_hd__nor2_1 _1330_ (.A(net43),
    .B(net38),
    .Y(_0671_));
 sky130_fd_sc_hd__a211oi_1 _1331_ (.A1(_0544_),
    .A2(_0548_),
    .B1(_0669_),
    .C1(_0671_),
    .Y(_0186_));
 sky130_fd_sc_hd__nand2_1 _1332_ (.A(\Dead_Time_Generator_inst_3.count_dt[1] ),
    .B(_0669_),
    .Y(_0672_));
 sky130_fd_sc_hd__or2_1 _1333_ (.A(\Dead_Time_Generator_inst_3.count_dt[1] ),
    .B(_0669_),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_1 _1334_ (.A(_0672_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__a21oi_1 _1335_ (.A1(_0545_),
    .A2(_0549_),
    .B1(_0674_),
    .Y(_0187_));
 sky130_fd_sc_hd__xnor2_1 _1336_ (.A(_0661_),
    .B(_0672_),
    .Y(_0675_));
 sky130_fd_sc_hd__a21oi_1 _1337_ (.A1(_0545_),
    .A2(_0549_),
    .B1(_0675_),
    .Y(_0188_));
 sky130_fd_sc_hd__and4_1 _1338_ (.A(\Dead_Time_Generator_inst_3.count_dt[3] ),
    .B(\Dead_Time_Generator_inst_3.count_dt[2] ),
    .C(\Dead_Time_Generator_inst_3.count_dt[1] ),
    .D(_0669_),
    .X(_0198_));
 sky130_fd_sc_hd__o21a_1 _1339_ (.A1(_0661_),
    .A2(_0672_),
    .B1(_0660_),
    .X(_0199_));
 sky130_fd_sc_hd__a211oi_1 _1340_ (.A1(_0544_),
    .A2(_0548_),
    .B1(_0198_),
    .C1(_0199_),
    .Y(_0189_));
 sky130_fd_sc_hd__o2bb2a_1 _1341_ (.A1_N(_0545_),
    .A2_N(_0549_),
    .B1(_0198_),
    .B2(net56),
    .X(_0190_));
 sky130_fd_sc_hd__and3_1 _1342_ (.A(_0625_),
    .B(_0626_),
    .C(_0645_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _1343_ (.A(_0200_),
    .X(_0191_));
 sky130_fd_sc_hd__and3_1 _1344_ (.A(\Dead_Time_Generator_inst_4.count_dt[0] ),
    .B(_0486_),
    .C(_0496_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _1345_ (.A(_0488_),
    .B(_0497_),
    .X(_0202_));
 sky130_fd_sc_hd__nor2_1 _1346_ (.A(_0201_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__and3_1 _1347_ (.A(_0545_),
    .B(_0549_),
    .C(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__clkbuf_1 _1348_ (.A(_0204_),
    .X(_0192_));
 sky130_fd_sc_hd__xor2_1 _1349_ (.A(\Dead_Time_Generator_inst_4.count_dt[1] ),
    .B(_0201_),
    .X(_0205_));
 sky130_fd_sc_hd__and3_1 _1350_ (.A(_0545_),
    .B(_0549_),
    .C(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _1351_ (.A(_0206_),
    .X(_0193_));
 sky130_fd_sc_hd__and3_1 _1352_ (.A(\Dead_Time_Generator_inst_4.count_dt[2] ),
    .B(\Dead_Time_Generator_inst_4.count_dt[1] ),
    .C(_0201_),
    .X(_0207_));
 sky130_fd_sc_hd__a21o_1 _1353_ (.A1(\Dead_Time_Generator_inst_4.count_dt[1] ),
    .A2(_0201_),
    .B1(\Dead_Time_Generator_inst_4.count_dt[2] ),
    .X(_0208_));
 sky130_fd_sc_hd__and2b_1 _1354_ (.A_N(_0207_),
    .B(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__and3_1 _1355_ (.A(_0545_),
    .B(_0549_),
    .C(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _1356_ (.A(_0210_),
    .X(_0194_));
 sky130_fd_sc_hd__xnor2_1 _1357_ (.A(_0487_),
    .B(_0207_),
    .Y(_0211_));
 sky130_fd_sc_hd__and3_1 _1358_ (.A(_0545_),
    .B(_0549_),
    .C(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _1359_ (.A(_0212_),
    .X(_0195_));
 sky130_fd_sc_hd__a21o_1 _1360_ (.A1(\Dead_Time_Generator_inst_4.count_dt[3] ),
    .A2(_0207_),
    .B1(\Dead_Time_Generator_inst_4.count_dt[4] ),
    .X(_0213_));
 sky130_fd_sc_hd__and3_1 _1361_ (.A(_0545_),
    .B(_0549_),
    .C(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _1362_ (.A(_0214_),
    .X(_0196_));
 sky130_fd_sc_hd__a21oi_1 _1363_ (.A1(_0545_),
    .A2(_0549_),
    .B1(net38),
    .Y(_0197_));
 sky130_fd_sc_hd__dfstp_1 _1364_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net34),
    .SET_B(_0064_),
    .Q(PMOS1_PS1_prev));
 sky130_fd_sc_hd__dfrtp_1 _1365_ (.CLK(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0002_),
    .RESET_B(_0065_),
    .Q(NMOS2_PS1_prev));
 sky130_fd_sc_hd__dfstp_1 _1366_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net32),
    .SET_B(_0066_),
    .Q(PMOS2_PS1_prev));
 sky130_fd_sc_hd__dfrtp_1 _1367_ (.CLK(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0000_),
    .RESET_B(_0067_),
    .Q(NMOS1_PS1_prev));
 sky130_fd_sc_hd__dfstp_1 _1368_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net84),
    .SET_B(_0068_),
    .Q(PMOS1_PS2_prev));
 sky130_fd_sc_hd__dfrtp_1 _1369_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0003_),
    .RESET_B(_0069_),
    .Q(NMOS2_PS2_prev));
 sky130_fd_sc_hd__dfstp_1 _1370_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0007_),
    .SET_B(_0070_),
    .Q(PMOS2_PS2_prev));
 sky130_fd_sc_hd__dfrtp_1 _1371_ (.CLK(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0001_),
    .RESET_B(_0071_),
    .Q(NMOS1_PS2_prev));
 sky130_fd_sc_hd__dfrtp_1 _1372_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0151_),
    .RESET_B(_0072_),
    .Q(\Shift_Register_Inst.data_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1373_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0152_),
    .RESET_B(_0073_),
    .Q(\Shift_Register_Inst.data_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1374_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0153_),
    .RESET_B(_0074_),
    .Q(\Shift_Register_Inst.data_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1375_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0154_),
    .RESET_B(_0075_),
    .Q(\Shift_Register_Inst.data_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1376_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0155_),
    .RESET_B(_0076_),
    .Q(\Shift_Register_Inst.data_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1377_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0156_),
    .RESET_B(_0077_),
    .Q(\Shift_Register_Inst.data_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1378_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0157_),
    .RESET_B(_0078_),
    .Q(\Shift_Register_Inst.data_out[11] ));
 sky130_fd_sc_hd__dfrtp_2 _1379_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0158_),
    .RESET_B(_0079_),
    .Q(\Shift_Register_Inst.data_out[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1380_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0159_),
    .RESET_B(_0080_),
    .Q(\Shift_Register_Inst.data_out[9] ));
 sky130_fd_sc_hd__dfrtp_4 _1381_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0160_),
    .RESET_B(_0081_),
    .Q(\Shift_Register_Inst.data_out[8] ));
 sky130_fd_sc_hd__dfrtp_2 _1382_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0161_),
    .RESET_B(_0082_),
    .Q(\Shift_Register_Inst.data_out[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1383_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0162_),
    .RESET_B(_0083_),
    .Q(\Shift_Register_Inst.data_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1384_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0163_),
    .RESET_B(_0084_),
    .Q(\Shift_Register_Inst.data_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1385_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0164_),
    .RESET_B(_0085_),
    .Q(\Dead_Time_Generator_inst_1.dt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1386_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0165_),
    .RESET_B(_0086_),
    .Q(\Dead_Time_Generator_inst_1.dt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1387_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0166_),
    .RESET_B(_0087_),
    .Q(\Dead_Time_Generator_inst_1.dt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1388_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0167_),
    .RESET_B(_0088_),
    .Q(\Dead_Time_Generator_inst_1.dt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1389_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0168_),
    .RESET_B(_0089_),
    .Q(\Shift_Register_Inst.shift_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1390_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0169_),
    .RESET_B(_0090_),
    .Q(\Shift_Register_Inst.shift_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1391_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0170_),
    .RESET_B(_0091_),
    .Q(\Shift_Register_Inst.shift_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1392_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0171_),
    .RESET_B(_0092_),
    .Q(\Shift_Register_Inst.shift_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1393_ (.CLK(clknet_1_1__leaf_CLK_SR),
    .D(_0172_),
    .RESET_B(_0093_),
    .Q(\Shift_Register_Inst.shift_state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1394_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0173_),
    .Q(\Dead_Time_Generator_inst_4.go ));
 sky130_fd_sc_hd__dfstp_2 _1395_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0014_),
    .SET_B(_0094_),
    .Q(\Signal_Generator_1_0phase_inst.direction ));
 sky130_fd_sc_hd__dfrtp_2 _1396_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0008_),
    .RESET_B(_0095_),
    .Q(\Signal_Generator_1_0phase_inst.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1397_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0009_),
    .RESET_B(_0096_),
    .Q(\Signal_Generator_1_0phase_inst.count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1398_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0010_),
    .RESET_B(_0097_),
    .Q(\Signal_Generator_1_0phase_inst.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1399_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0011_),
    .RESET_B(_0098_),
    .Q(\Signal_Generator_1_0phase_inst.count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1400_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0012_),
    .RESET_B(_0099_),
    .Q(\Signal_Generator_1_0phase_inst.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1401_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0013_),
    .RESET_B(_0100_),
    .Q(\Signal_Generator_1_0phase_inst.count[5] ));
 sky130_fd_sc_hd__dfstp_1 _1402_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0035_),
    .SET_B(_0101_),
    .Q(\Signal_Generator_1_90phase_inst.direction ));
 sky130_fd_sc_hd__dfstp_1 _1403_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0029_),
    .SET_B(_0102_),
    .Q(\Signal_Generator_1_90phase_inst.count[0] ));
 sky130_fd_sc_hd__dfstp_1 _1404_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0030_),
    .SET_B(_0103_),
    .Q(\Signal_Generator_1_90phase_inst.count[1] ));
 sky130_fd_sc_hd__dfstp_2 _1405_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0031_),
    .SET_B(_0104_),
    .Q(\Signal_Generator_1_90phase_inst.count[2] ));
 sky130_fd_sc_hd__dfstp_1 _1406_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0032_),
    .SET_B(_0105_),
    .Q(\Signal_Generator_1_90phase_inst.count[3] ));
 sky130_fd_sc_hd__dfstp_2 _1407_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0033_),
    .SET_B(_0106_),
    .Q(\Signal_Generator_1_90phase_inst.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1408_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0034_),
    .RESET_B(_0107_),
    .Q(\Signal_Generator_1_90phase_inst.count[5] ));
 sky130_fd_sc_hd__dfstp_1 _1409_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0021_),
    .SET_B(_0108_),
    .Q(\Signal_Generator_1_180phase_inst.direction ));
 sky130_fd_sc_hd__dfstp_1 _1410_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0015_),
    .SET_B(_0109_),
    .Q(\Signal_Generator_1_180phase_inst.count[0] ));
 sky130_fd_sc_hd__dfstp_1 _1411_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0016_),
    .SET_B(_0110_),
    .Q(\Signal_Generator_1_180phase_inst.count[1] ));
 sky130_fd_sc_hd__dfstp_2 _1412_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0017_),
    .SET_B(_0111_),
    .Q(\Signal_Generator_1_180phase_inst.count[2] ));
 sky130_fd_sc_hd__dfstp_1 _1413_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0018_),
    .SET_B(_0112_),
    .Q(\Signal_Generator_1_180phase_inst.count[3] ));
 sky130_fd_sc_hd__dfstp_2 _1414_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0019_),
    .SET_B(_0113_),
    .Q(\Signal_Generator_1_180phase_inst.count[4] ));
 sky130_fd_sc_hd__dfstp_1 _1415_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0020_),
    .SET_B(_0114_),
    .Q(\Signal_Generator_1_180phase_inst.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1416_ (.CLK(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0028_),
    .RESET_B(_0115_),
    .Q(\Signal_Generator_1_270phase_inst.direction ));
 sky130_fd_sc_hd__dfrtp_2 _1417_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0022_),
    .RESET_B(_0116_),
    .Q(\Signal_Generator_1_270phase_inst.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1418_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0023_),
    .RESET_B(_0117_),
    .Q(\Signal_Generator_1_270phase_inst.count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1419_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0024_),
    .RESET_B(_0118_),
    .Q(\Signal_Generator_1_270phase_inst.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1420_ (.CLK(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0025_),
    .RESET_B(_0119_),
    .Q(\Signal_Generator_1_270phase_inst.count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1421_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0026_),
    .RESET_B(_0120_),
    .Q(\Signal_Generator_1_270phase_inst.count[4] ));
 sky130_fd_sc_hd__dfstp_1 _1422_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net78),
    .SET_B(_0121_),
    .Q(\Signal_Generator_1_270phase_inst.count[5] ));
 sky130_fd_sc_hd__dfstp_1 _1423_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0042_),
    .SET_B(_0122_),
    .Q(\Signal_Generator_2_0phase_inst.direction ));
 sky130_fd_sc_hd__dfrtp_2 _1424_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0036_),
    .RESET_B(_0123_),
    .Q(\Signal_Generator_2_0phase_inst.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1425_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0037_),
    .RESET_B(_0124_),
    .Q(\Signal_Generator_2_0phase_inst.count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1426_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0038_),
    .RESET_B(_0125_),
    .Q(\Signal_Generator_2_0phase_inst.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1427_ (.CLK(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0039_),
    .RESET_B(_0126_),
    .Q(\Signal_Generator_2_0phase_inst.count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1428_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0040_),
    .RESET_B(_0127_),
    .Q(\Signal_Generator_2_0phase_inst.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1429_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0041_),
    .RESET_B(_0128_),
    .Q(\Signal_Generator_2_0phase_inst.count[5] ));
 sky130_fd_sc_hd__dfstp_1 _1430_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0063_),
    .SET_B(_0129_),
    .Q(\Signal_Generator_2_90phase_inst.direction ));
 sky130_fd_sc_hd__dfstp_2 _1431_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0057_),
    .SET_B(_0130_),
    .Q(\Signal_Generator_2_90phase_inst.count[0] ));
 sky130_fd_sc_hd__dfstp_1 _1432_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0058_),
    .SET_B(_0131_),
    .Q(\Signal_Generator_2_90phase_inst.count[1] ));
 sky130_fd_sc_hd__dfstp_2 _1433_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0059_),
    .SET_B(_0132_),
    .Q(\Signal_Generator_2_90phase_inst.count[2] ));
 sky130_fd_sc_hd__dfstp_1 _1434_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0060_),
    .SET_B(_0133_),
    .Q(\Signal_Generator_2_90phase_inst.count[3] ));
 sky130_fd_sc_hd__dfstp_2 _1435_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0061_),
    .SET_B(_0134_),
    .Q(\Signal_Generator_2_90phase_inst.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1436_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0062_),
    .RESET_B(_0135_),
    .Q(\Signal_Generator_2_90phase_inst.count[5] ));
 sky130_fd_sc_hd__dfstp_1 _1437_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0049_),
    .SET_B(_0136_),
    .Q(\Signal_Generator_2_180phase_inst.direction ));
 sky130_fd_sc_hd__dfstp_1 _1438_ (.CLK(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0043_),
    .SET_B(_0137_),
    .Q(\Signal_Generator_2_180phase_inst.count[0] ));
 sky130_fd_sc_hd__dfstp_1 _1439_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0044_),
    .SET_B(_0138_),
    .Q(\Signal_Generator_2_180phase_inst.count[1] ));
 sky130_fd_sc_hd__dfstp_2 _1440_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0045_),
    .SET_B(_0139_),
    .Q(\Signal_Generator_2_180phase_inst.count[2] ));
 sky130_fd_sc_hd__dfstp_1 _1441_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0046_),
    .SET_B(_0140_),
    .Q(\Signal_Generator_2_180phase_inst.count[3] ));
 sky130_fd_sc_hd__dfstp_2 _1442_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0047_),
    .SET_B(_0141_),
    .Q(\Signal_Generator_2_180phase_inst.count[4] ));
 sky130_fd_sc_hd__dfstp_1 _1443_ (.CLK(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0048_),
    .SET_B(_0142_),
    .Q(\Signal_Generator_2_180phase_inst.count[5] ));
 sky130_fd_sc_hd__dfrtp_4 _1444_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0056_),
    .RESET_B(_0143_),
    .Q(\Signal_Generator_2_270phase_inst.direction ));
 sky130_fd_sc_hd__dfrtp_2 _1445_ (.CLK(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0050_),
    .RESET_B(_0144_),
    .Q(\Signal_Generator_2_270phase_inst.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1446_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0051_),
    .RESET_B(_0145_),
    .Q(\Signal_Generator_2_270phase_inst.count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1447_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0052_),
    .RESET_B(_0146_),
    .Q(\Signal_Generator_2_270phase_inst.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1448_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0053_),
    .RESET_B(_0147_),
    .Q(\Signal_Generator_2_270phase_inst.count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1449_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0054_),
    .RESET_B(_0148_),
    .Q(\Signal_Generator_2_270phase_inst.count[4] ));
 sky130_fd_sc_hd__dfstp_1 _1450_ (.CLK(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0055_),
    .SET_B(_0149_),
    .Q(\Signal_Generator_2_270phase_inst.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1451_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net42),
    .Q(\Dead_Time_Generator_inst_1.count_dt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1452_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0175_),
    .Q(\Dead_Time_Generator_inst_1.count_dt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1453_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0176_),
    .Q(\Dead_Time_Generator_inst_1.count_dt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1454_ (.CLK(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net55),
    .Q(\Dead_Time_Generator_inst_1.count_dt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1455_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0178_),
    .Q(\Dead_Time_Generator_inst_1.count_dt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1456_ (.CLK(clknet_1_0__leaf_CLK_SR),
    .D(_0179_),
    .RESET_B(_0150_),
    .Q(\Dead_Time_Generator_inst_1.dt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1457_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0180_),
    .Q(\Dead_Time_Generator_inst_2.count_dt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1458_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0181_),
    .Q(\Dead_Time_Generator_inst_2.count_dt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1459_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0182_),
    .Q(\Dead_Time_Generator_inst_2.count_dt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1460_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0183_),
    .Q(\Dead_Time_Generator_inst_2.count_dt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1461_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0184_),
    .Q(\Dead_Time_Generator_inst_2.count_dt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1462_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0185_),
    .Q(\Dead_Time_Generator_inst_1.go ));
 sky130_fd_sc_hd__dfxtp_1 _1463_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net44),
    .Q(\Dead_Time_Generator_inst_3.count_dt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1464_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0187_),
    .Q(\Dead_Time_Generator_inst_3.count_dt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1465_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0188_),
    .Q(\Dead_Time_Generator_inst_3.count_dt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1466_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(net72),
    .Q(\Dead_Time_Generator_inst_3.count_dt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1467_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0190_),
    .Q(\Dead_Time_Generator_inst_3.count_dt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1468_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0191_),
    .Q(\Dead_Time_Generator_inst_2.go ));
 sky130_fd_sc_hd__dfxtp_1 _1469_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0192_),
    .Q(\Dead_Time_Generator_inst_4.count_dt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1470_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0193_),
    .Q(\Dead_Time_Generator_inst_4.count_dt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1471_ (.CLK(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0194_),
    .Q(\Dead_Time_Generator_inst_4.count_dt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1472_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0195_),
    .Q(\Dead_Time_Generator_inst_4.count_dt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1473_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0196_),
    .Q(\Dead_Time_Generator_inst_4.count_dt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1474_ (.CLK(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ),
    .D(_0197_),
    .Q(\Dead_Time_Generator_inst_3.go ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK_SR (.A(CLK_SR),
    .X(clknet_0_CLK_SR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_Dead_Time_Generator_inst_1.clk  (.A(\Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_0_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_CLK_SR (.A(clknet_0_CLK_SR),
    .X(clknet_1_0__leaf_CLK_SR));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_CLK_SR (.A(clknet_0_CLK_SR),
    .X(clknet_1_1__leaf_CLK_SR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_Dead_Time_Generator_inst_1.clk  (.A(\clknet_0_Dead_Time_Generator_inst_1.clk ),
    .X(\clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk ));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\Dead_Time_Generator_inst_3.go ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\Dead_Time_Generator_inst_1.go ),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 hold12 (.A(net86),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0670_),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 hold14 (.A(\Dead_Time_Generator_inst_1.dt[3] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0621_),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\Shift_Register_Inst.data_out[16] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0174_),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\Dead_Time_Generator_inst_3.count_dt[0] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0186_),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\Dead_Time_Generator_inst_1.dt[3] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0494_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0496_),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\Signal_Generator_1_270phase_inst.count[0] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\Signal_Generator_2_270phase_inst.count[0] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\Dead_Time_Generator_inst_1.count_dt[4] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\Signal_Generator_2_90phase_inst.count[0] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\Signal_Generator_1_0phase_inst.count[0] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\Dead_Time_Generator_inst_1.dt[4] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\Dead_Time_Generator_inst_1.count_dt[3] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0177_),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\Dead_Time_Generator_inst_3.count_dt[4] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\Signal_Generator_2_180phase_inst.count[0] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\Signal_Generator_2_0phase_inst.count[0] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\Signal_Generator_1_180phase_inst.count[0] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\Signal_Generator_1_90phase_inst.count[0] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\Shift_Register_Inst.shift_state[4] ),
    .X(net61));
 sky130_fd_sc_hd__buf_1 hold37 (.A(\Signal_Generator_2_180phase_inst.direction ),
    .X(net62));
 sky130_fd_sc_hd__buf_1 hold38 (.A(\Signal_Generator_1_90phase_inst.direction ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\Shift_Register_Inst.shift_state[1] ),
    .X(net64));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold40 (.A(\Signal_Generator_2_90phase_inst.direction ),
    .X(net65));
 sky130_fd_sc_hd__buf_1 hold41 (.A(\Signal_Generator_1_180phase_inst.direction ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\Shift_Register_Inst.shift_state[0] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\Signal_Generator_1_270phase_inst.direction ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\Signal_Generator_2_0phase_inst.direction ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\Dead_Time_Generator_inst_1.count_dt[2] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\Dead_Time_Generator_inst_3.count_dt[3] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0189_),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\Signal_Generator_1_0phase_inst.count[4] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\Dead_Time_Generator_inst_3.count_dt[2] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\Shift_Register_Inst.data_out[15] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\Signal_Generator_1_0phase_inst.direction ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\Shift_Register_Inst.data_out[14] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\Signal_Generator_1_270phase_inst.direction ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0027_),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\Shift_Register_Inst.data_out[15] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\Signal_Generator_2_0phase_inst.direction ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\Signal_Generator_2_90phase_inst.direction ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\Signal_Generator_1_180phase_inst.direction ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\Signal_Generator_2_180phase_inst.direction ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0005_),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold6 (.A(net30),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\Shift_Register_Inst.data_out[13] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\Dead_Time_Generator_inst_1.dt[4] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0006_),
    .X(net32));
 sky130_fd_sc_hd__buf_1 hold8 (.A(net85),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0004_),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input1 (.A(Data_SR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(d2[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(d2[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(d2[3]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(d2[4]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(d2[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(RST),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(d1[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(d1[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(d1[2]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(d1[3]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(d1[4]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(d1[5]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(d2[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(NMOS1_PS1));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(NMOS1_PS2));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(NMOS2_PS1));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(NMOS2_PS2));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(NMOS_PS3));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(PMOS1_PS1));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(PMOS1_PS2));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(PMOS2_PS1));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(PMOS2_PS2));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(PMOS_PS3));
 sky130_fd_sc_hd__buf_6 output25 (.A(net25),
    .X(SIGNAL_OUTPUT));
endmodule

