magic
tech sky130A
magscale 1 2
timestamp 1697513884
<< viali >>
rect 3985 27081 4019 27115
rect 7389 27081 7423 27115
rect 12081 27081 12115 27115
rect 19625 27081 19659 27115
rect 23489 27081 23523 27115
rect 3893 27013 3927 27047
rect 1409 26945 1443 26979
rect 7297 26945 7331 26979
rect 11897 26945 11931 26979
rect 15761 26945 15795 26979
rect 19533 26945 19567 26979
rect 23397 26945 23431 26979
rect 1593 26741 1627 26775
rect 15577 26741 15611 26775
rect 9689 26469 9723 26503
rect 6837 26401 6871 26435
rect 16313 26401 16347 26435
rect 17325 26401 17359 26435
rect 17509 26401 17543 26435
rect 20269 26401 20303 26435
rect 6561 26333 6595 26367
rect 9965 26333 9999 26367
rect 12081 26333 12115 26367
rect 12449 26333 12483 26367
rect 15301 26333 15335 26367
rect 15761 26333 15795 26367
rect 17233 26333 17267 26367
rect 17417 26333 17451 26367
rect 18061 26333 18095 26367
rect 20177 26333 20211 26367
rect 20453 26333 20487 26367
rect 9229 26265 9263 26299
rect 9413 26265 9447 26299
rect 9689 26265 9723 26299
rect 9873 26265 9907 26299
rect 15393 26265 15427 26299
rect 17693 26265 17727 26299
rect 17877 26265 17911 26299
rect 20545 26265 20579 26299
rect 8309 26197 8343 26231
rect 9597 26197 9631 26231
rect 13875 26197 13909 26231
rect 17049 26197 17083 26231
rect 9689 25993 9723 26027
rect 13829 25993 13863 26027
rect 21925 25993 21959 26027
rect 6653 25925 6687 25959
rect 9321 25925 9355 25959
rect 19073 25925 19107 25959
rect 6377 25857 6411 25891
rect 8677 25857 8711 25891
rect 9137 25857 9171 25891
rect 9413 25857 9447 25891
rect 9505 25857 9539 25891
rect 9965 25857 9999 25891
rect 10425 25857 10459 25891
rect 10609 25857 10643 25891
rect 11529 25857 11563 25891
rect 11805 25857 11839 25891
rect 13737 25857 13771 25891
rect 16313 25857 16347 25891
rect 16773 25857 16807 25891
rect 17417 25857 17451 25891
rect 18981 25857 19015 25891
rect 19717 25857 19751 25891
rect 22109 25857 22143 25891
rect 22201 25857 22235 25891
rect 8401 25789 8435 25823
rect 8769 25789 8803 25823
rect 9045 25789 9079 25823
rect 9873 25789 9907 25823
rect 12173 25789 12207 25823
rect 14381 25789 14415 25823
rect 14749 25789 14783 25823
rect 17049 25789 17083 25823
rect 20085 25789 20119 25823
rect 22569 25789 22603 25823
rect 10333 25721 10367 25755
rect 16405 25721 16439 25755
rect 10425 25653 10459 25687
rect 11621 25653 11655 25687
rect 13553 25653 13587 25687
rect 16175 25653 16209 25687
rect 16865 25653 16899 25687
rect 18797 25653 18831 25687
rect 21465 25653 21499 25687
rect 23995 25653 24029 25687
rect 6929 25449 6963 25483
rect 7481 25449 7515 25483
rect 9781 25449 9815 25483
rect 12725 25449 12759 25483
rect 15485 25449 15519 25483
rect 23673 25449 23707 25483
rect 9137 25381 9171 25415
rect 9873 25381 9907 25415
rect 13277 25381 13311 25415
rect 13553 25381 13587 25415
rect 23029 25381 23063 25415
rect 4721 25313 4755 25347
rect 10517 25313 10551 25347
rect 12265 25313 12299 25347
rect 15577 25313 15611 25347
rect 16773 25313 16807 25347
rect 17141 25313 17175 25347
rect 19441 25313 19475 25347
rect 21373 25313 21407 25347
rect 6837 25245 6871 25279
rect 7389 25245 7423 25279
rect 9137 25245 9171 25279
rect 9321 25245 9355 25279
rect 9597 25245 9631 25279
rect 9873 25245 9907 25279
rect 10057 25245 10091 25279
rect 10149 25245 10183 25279
rect 10241 25245 10275 25279
rect 12633 25245 12667 25279
rect 13277 25245 13311 25279
rect 13461 25245 13495 25279
rect 13829 25245 13863 25279
rect 14565 25245 14599 25279
rect 14933 25245 14967 25279
rect 15117 25245 15151 25279
rect 15301 25245 15335 25279
rect 15761 25245 15795 25279
rect 16037 25245 16071 25279
rect 16681 25245 16715 25279
rect 17509 25245 17543 25279
rect 21465 25245 21499 25279
rect 22477 25245 22511 25279
rect 23305 25245 23339 25279
rect 23581 25245 23615 25279
rect 24409 25245 24443 25279
rect 25789 25245 25823 25279
rect 4997 25177 5031 25211
rect 6745 25177 6779 25211
rect 9413 25177 9447 25211
rect 13553 25177 13587 25211
rect 15209 25177 15243 25211
rect 19717 25177 19751 25211
rect 23121 25177 23155 25211
rect 13737 25109 13771 25143
rect 14749 25109 14783 25143
rect 15945 25109 15979 25143
rect 17049 25109 17083 25143
rect 18935 25109 18969 25143
rect 21189 25109 21223 25143
rect 21833 25109 21867 25143
rect 23489 25109 23523 25143
rect 25053 25109 25087 25143
rect 25973 25109 26007 25143
rect 7113 24905 7147 24939
rect 9429 24905 9463 24939
rect 13093 24905 13127 24939
rect 14013 24905 14047 24939
rect 15485 24905 15519 24939
rect 16497 24905 16531 24939
rect 16957 24905 16991 24939
rect 17785 24905 17819 24939
rect 19717 24905 19751 24939
rect 20361 24905 20395 24939
rect 9229 24837 9263 24871
rect 12909 24837 12943 24871
rect 14381 24837 14415 24871
rect 16129 24837 16163 24871
rect 16345 24837 16379 24871
rect 17443 24837 17477 24871
rect 20729 24837 20763 24871
rect 5825 24769 5859 24803
rect 5917 24769 5951 24803
rect 6745 24769 6779 24803
rect 7389 24769 7423 24803
rect 7573 24769 7607 24803
rect 7665 24769 7699 24803
rect 7849 24769 7883 24803
rect 8033 24769 8067 24803
rect 8401 24769 8435 24803
rect 8953 24769 8987 24803
rect 9873 24769 9907 24803
rect 13185 24769 13219 24803
rect 13645 24769 13679 24803
rect 13829 24769 13863 24803
rect 14105 24769 14139 24803
rect 14289 24769 14323 24803
rect 14473 24769 14507 24803
rect 14749 24769 14783 24803
rect 14933 24769 14967 24803
rect 15393 24769 15427 24803
rect 15577 24769 15611 24803
rect 16681 24769 16715 24803
rect 16773 24769 16807 24803
rect 17141 24769 17175 24803
rect 17233 24769 17267 24803
rect 17325 24769 17359 24803
rect 17969 24769 18003 24803
rect 18061 24769 18095 24803
rect 18245 24769 18279 24803
rect 18429 24769 18463 24803
rect 18613 24769 18647 24803
rect 18705 24769 18739 24803
rect 18889 24769 18923 24803
rect 19073 24769 19107 24803
rect 19165 24769 19199 24803
rect 19993 24769 20027 24803
rect 20545 24769 20579 24803
rect 20637 24769 20671 24803
rect 20847 24769 20881 24803
rect 21005 24769 21039 24803
rect 21281 24769 21315 24803
rect 21557 24769 21591 24803
rect 22109 24769 22143 24803
rect 22201 24769 22235 24803
rect 22385 24769 22419 24803
rect 22569 24769 22603 24803
rect 6837 24701 6871 24735
rect 9689 24701 9723 24735
rect 10057 24701 10091 24735
rect 15117 24701 15151 24735
rect 17601 24701 17635 24735
rect 19901 24701 19935 24735
rect 20085 24701 20119 24735
rect 20177 24701 20211 24735
rect 22661 24701 22695 24735
rect 7481 24633 7515 24667
rect 14657 24633 14691 24667
rect 18153 24633 18187 24667
rect 18797 24633 18831 24667
rect 21373 24633 21407 24667
rect 21465 24633 21499 24667
rect 22293 24633 22327 24667
rect 7205 24565 7239 24599
rect 8217 24565 8251 24599
rect 8493 24565 8527 24599
rect 9045 24565 9079 24599
rect 9413 24565 9447 24599
rect 9597 24565 9631 24599
rect 12909 24565 12943 24599
rect 16313 24565 16347 24599
rect 21097 24565 21131 24599
rect 21925 24565 21959 24599
rect 7573 24361 7607 24395
rect 8585 24361 8619 24395
rect 8769 24361 8803 24395
rect 14657 24361 14691 24395
rect 15025 24361 15059 24395
rect 15117 24361 15151 24395
rect 15577 24361 15611 24395
rect 15761 24361 15795 24395
rect 15945 24361 15979 24395
rect 17325 24361 17359 24395
rect 20637 24361 20671 24395
rect 21097 24361 21131 24395
rect 22477 24361 22511 24395
rect 13875 24293 13909 24327
rect 17785 24293 17819 24327
rect 23765 24293 23799 24327
rect 5641 24225 5675 24259
rect 10241 24225 10275 24259
rect 12449 24225 12483 24259
rect 14197 24225 14231 24259
rect 14887 24225 14921 24259
rect 15485 24225 15519 24259
rect 16221 24225 16255 24259
rect 16405 24225 16439 24259
rect 17509 24225 17543 24259
rect 20821 24225 20855 24259
rect 21281 24225 21315 24259
rect 6009 24157 6043 24191
rect 7774 24167 7808 24201
rect 7941 24157 7975 24191
rect 8217 24157 8251 24191
rect 9137 24157 9171 24191
rect 9413 24157 9447 24191
rect 9505 24157 9539 24191
rect 9781 24157 9815 24191
rect 9873 24157 9907 24191
rect 12081 24157 12115 24191
rect 14289 24157 14323 24191
rect 14749 24157 14783 24191
rect 15209 24157 15243 24191
rect 15577 24157 15611 24191
rect 16129 24157 16163 24191
rect 16313 24157 16347 24191
rect 17233 24157 17267 24191
rect 20545 24157 20579 24191
rect 21189 24157 21223 24191
rect 22477 24157 22511 24191
rect 22661 24157 22695 24191
rect 23121 24157 23155 24191
rect 23489 24157 23523 24191
rect 23949 24157 23983 24191
rect 24041 24157 24075 24191
rect 24409 24157 24443 24191
rect 7849 24089 7883 24123
rect 8079 24089 8113 24123
rect 8401 24089 8435 24123
rect 8953 24089 8987 24123
rect 9689 24089 9723 24123
rect 10517 24089 10551 24123
rect 15301 24089 15335 24123
rect 23305 24089 23339 24123
rect 23397 24089 23431 24123
rect 23765 24089 23799 24123
rect 7435 24021 7469 24055
rect 8601 24021 8635 24055
rect 9321 24021 9355 24055
rect 10057 24021 10091 24055
rect 11989 24021 12023 24055
rect 23673 24021 23707 24055
rect 24501 24021 24535 24055
rect 6561 23817 6595 23851
rect 6837 23817 6871 23851
rect 8309 23817 8343 23851
rect 8493 23817 8527 23851
rect 10425 23817 10459 23851
rect 11621 23817 11655 23851
rect 13093 23817 13127 23851
rect 15025 23817 15059 23851
rect 15777 23817 15811 23851
rect 15945 23817 15979 23851
rect 20913 23817 20947 23851
rect 22385 23817 22419 23851
rect 22937 23817 22971 23851
rect 4261 23749 4295 23783
rect 4445 23749 4479 23783
rect 5181 23749 5215 23783
rect 9806 23749 9840 23783
rect 15577 23749 15611 23783
rect 21097 23749 21131 23783
rect 21313 23749 21347 23783
rect 22753 23749 22787 23783
rect 5365 23681 5399 23715
rect 6469 23681 6503 23715
rect 7021 23681 7055 23715
rect 7297 23681 7331 23715
rect 7757 23681 7791 23715
rect 8125 23681 8159 23715
rect 8677 23681 8711 23715
rect 8861 23681 8895 23715
rect 8953 23681 8987 23715
rect 9229 23681 9263 23715
rect 9689 23687 9723 23721
rect 9965 23681 9999 23715
rect 10057 23681 10091 23715
rect 11529 23681 11563 23715
rect 13001 23681 13035 23715
rect 13829 23681 13863 23715
rect 14289 23681 14323 23715
rect 14473 23681 14507 23715
rect 14749 23681 14783 23715
rect 14841 23681 14875 23715
rect 20729 23681 20763 23715
rect 21005 23681 21039 23715
rect 22201 23681 22235 23715
rect 22477 23681 22511 23715
rect 22569 23681 22603 23715
rect 23397 23681 23431 23715
rect 4169 23613 4203 23647
rect 7113 23613 7147 23647
rect 7205 23613 7239 23647
rect 9367 23613 9401 23647
rect 9597 23613 9631 23647
rect 10609 23613 10643 23647
rect 10701 23613 10735 23647
rect 10793 23613 10827 23647
rect 10885 23613 10919 23647
rect 13921 23613 13955 23647
rect 14381 23613 14415 23647
rect 23029 23613 23063 23647
rect 4721 23545 4755 23579
rect 5549 23545 5583 23579
rect 8773 23545 8807 23579
rect 9505 23545 9539 23579
rect 14197 23545 14231 23579
rect 21465 23545 21499 23579
rect 3709 23477 3743 23511
rect 8125 23477 8159 23511
rect 9965 23477 9999 23511
rect 10241 23477 10275 23511
rect 15761 23477 15795 23511
rect 20545 23477 20579 23511
rect 21281 23477 21315 23511
rect 22201 23477 22235 23511
rect 24777 23477 24811 23511
rect 5549 23273 5583 23307
rect 9873 23273 9907 23307
rect 17141 23273 17175 23307
rect 20821 23273 20855 23307
rect 20913 23273 20947 23307
rect 21741 23273 21775 23307
rect 22661 23273 22695 23307
rect 23121 23273 23155 23307
rect 23765 23273 23799 23307
rect 21925 23205 21959 23239
rect 5641 23137 5675 23171
rect 20085 23137 20119 23171
rect 21189 23137 21223 23171
rect 21281 23137 21315 23171
rect 22201 23137 22235 23171
rect 23489 23137 23523 23171
rect 23949 23137 23983 23171
rect 3801 23069 3835 23103
rect 6377 23069 6411 23103
rect 9781 23069 9815 23103
rect 9965 23069 9999 23103
rect 16773 23069 16807 23103
rect 18153 23069 18187 23103
rect 18337 23069 18371 23103
rect 18429 23069 18463 23103
rect 19993 23069 20027 23103
rect 20177 23069 20211 23103
rect 20315 23069 20349 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 21097 23069 21131 23103
rect 21373 23069 21407 23103
rect 22293 23069 22327 23103
rect 22937 23069 22971 23103
rect 23397 23069 23431 23103
rect 23857 23069 23891 23103
rect 24041 23069 24075 23103
rect 4077 23001 4111 23035
rect 6469 23001 6503 23035
rect 20545 23001 20579 23035
rect 21557 23001 21591 23035
rect 21773 23001 21807 23035
rect 22753 23001 22787 23035
rect 6285 22933 6319 22967
rect 17141 22933 17175 22967
rect 17325 22933 17359 22967
rect 17969 22933 18003 22967
rect 4077 22729 4111 22763
rect 4997 22729 5031 22763
rect 9965 22729 9999 22763
rect 11177 22729 11211 22763
rect 11729 22729 11763 22763
rect 11897 22729 11931 22763
rect 12465 22729 12499 22763
rect 13661 22729 13695 22763
rect 13829 22729 13863 22763
rect 18337 22729 18371 22763
rect 19717 22729 19751 22763
rect 22569 22729 22603 22763
rect 6009 22661 6043 22695
rect 9597 22661 9631 22695
rect 9797 22661 9831 22695
rect 10977 22661 11011 22695
rect 11529 22661 11563 22695
rect 12265 22661 12299 22695
rect 13461 22661 13495 22695
rect 15577 22661 15611 22695
rect 16221 22661 16255 22695
rect 17049 22661 17083 22695
rect 18889 22661 18923 22695
rect 24455 22661 24489 22695
rect 4261 22593 4295 22627
rect 4905 22593 4939 22627
rect 5733 22593 5767 22627
rect 10241 22593 10275 22627
rect 10517 22593 10551 22627
rect 15853 22593 15887 22627
rect 17417 22593 17451 22627
rect 18061 22593 18095 22627
rect 18153 22593 18187 22627
rect 18429 22593 18463 22627
rect 19257 22593 19291 22627
rect 19395 22593 19429 22627
rect 19717 22593 19751 22627
rect 22385 22593 22419 22627
rect 22661 22593 22695 22627
rect 23029 22593 23063 22627
rect 5181 22525 5215 22559
rect 12817 22525 12851 22559
rect 16681 22525 16715 22559
rect 17969 22525 18003 22559
rect 19809 22525 19843 22559
rect 20177 22525 20211 22559
rect 22201 22525 22235 22559
rect 4537 22457 4571 22491
rect 12633 22457 12667 22491
rect 15209 22457 15243 22491
rect 16405 22457 16439 22491
rect 17509 22457 17543 22491
rect 18521 22457 18555 22491
rect 19073 22457 19107 22491
rect 21603 22457 21637 22491
rect 9781 22389 9815 22423
rect 10333 22389 10367 22423
rect 10609 22389 10643 22423
rect 11161 22389 11195 22423
rect 11345 22389 11379 22423
rect 11713 22389 11747 22423
rect 12449 22389 12483 22423
rect 13369 22389 13403 22423
rect 13645 22389 13679 22423
rect 15577 22389 15611 22423
rect 15761 22389 15795 22423
rect 16221 22389 16255 22423
rect 17049 22389 17083 22423
rect 17233 22389 17267 22423
rect 17693 22389 17727 22423
rect 18889 22389 18923 22423
rect 19533 22389 19567 22423
rect 15945 22185 15979 22219
rect 16497 22185 16531 22219
rect 17601 22185 17635 22219
rect 17693 22185 17727 22219
rect 18521 22185 18555 22219
rect 18797 22185 18831 22219
rect 19717 22185 19751 22219
rect 20177 22185 20211 22219
rect 11161 22117 11195 22151
rect 17509 22117 17543 22151
rect 18337 22117 18371 22151
rect 5825 22049 5859 22083
rect 13829 22049 13863 22083
rect 15761 22049 15795 22083
rect 16313 22049 16347 22083
rect 18061 22049 18095 22083
rect 19809 22049 19843 22083
rect 21557 22049 21591 22083
rect 23765 22049 23799 22083
rect 3801 21981 3835 22015
rect 5733 21981 5767 22015
rect 5917 21981 5951 22015
rect 6009 21981 6043 22015
rect 6193 21981 6227 22015
rect 6929 21981 6963 22015
rect 8769 21981 8803 22015
rect 9137 21981 9171 22015
rect 9413 21981 9447 22015
rect 11437 21981 11471 22015
rect 11713 21981 11747 22015
rect 12081 21981 12115 22015
rect 14105 21981 14139 22015
rect 14473 21981 14507 22015
rect 15117 21981 15151 22015
rect 15209 21981 15243 22015
rect 15945 21981 15979 22015
rect 16221 21981 16255 22015
rect 16497 21981 16531 22015
rect 16865 21981 16899 22015
rect 17049 21981 17083 22015
rect 17785 21981 17819 22015
rect 17969 21981 18003 22015
rect 19993 21981 20027 22015
rect 21465 21981 21499 22015
rect 23673 21981 23707 22015
rect 9689 21913 9723 21947
rect 11529 21913 11563 21947
rect 12357 21913 12391 21947
rect 15669 21913 15703 21947
rect 16957 21913 16991 21947
rect 18613 21913 18647 21947
rect 18829 21913 18863 21947
rect 19717 21913 19751 21947
rect 3985 21845 4019 21879
rect 6193 21845 6227 21879
rect 7021 21845 7055 21879
rect 8585 21845 8619 21879
rect 8953 21845 8987 21879
rect 11897 21845 11931 21879
rect 14289 21845 14323 21879
rect 15301 21845 15335 21879
rect 16129 21845 16163 21879
rect 16681 21845 16715 21879
rect 17233 21845 17267 21879
rect 18981 21845 19015 21879
rect 8401 21641 8435 21675
rect 17693 21641 17727 21675
rect 6653 21573 6687 21607
rect 9597 21573 9631 21607
rect 11345 21573 11379 21607
rect 17509 21573 17543 21607
rect 3617 21505 3651 21539
rect 8769 21505 8803 21539
rect 8861 21505 8895 21539
rect 12449 21505 12483 21539
rect 14565 21505 14599 21539
rect 15301 21505 15335 21539
rect 15577 21505 15611 21539
rect 18153 21505 18187 21539
rect 18337 21505 18371 21539
rect 18613 21505 18647 21539
rect 25789 21505 25823 21539
rect 1501 21437 1535 21471
rect 1777 21437 1811 21471
rect 3525 21437 3559 21471
rect 3893 21437 3927 21471
rect 5365 21437 5399 21471
rect 5549 21437 5583 21471
rect 6377 21437 6411 21471
rect 8953 21437 8987 21471
rect 9321 21437 9355 21471
rect 12817 21437 12851 21471
rect 14381 21437 14415 21471
rect 15418 21437 15452 21471
rect 17141 21437 17175 21471
rect 18429 21437 18463 21471
rect 6193 21369 6227 21403
rect 14243 21369 14277 21403
rect 15025 21369 15059 21403
rect 18245 21369 18279 21403
rect 8125 21301 8159 21335
rect 16221 21301 16255 21335
rect 17509 21301 17543 21335
rect 17969 21301 18003 21335
rect 25973 21301 26007 21335
rect 2145 21097 2179 21131
rect 2513 21097 2547 21131
rect 3525 21097 3559 21131
rect 3801 21097 3835 21131
rect 4905 21097 4939 21131
rect 5089 21097 5123 21131
rect 7573 21097 7607 21131
rect 8033 21097 8067 21131
rect 8953 21097 8987 21131
rect 11897 21097 11931 21131
rect 13093 21097 13127 21131
rect 14381 21097 14415 21131
rect 16405 21097 16439 21131
rect 17877 21097 17911 21131
rect 21373 21097 21407 21131
rect 4537 21029 4571 21063
rect 7389 21029 7423 21063
rect 1961 20961 1995 20995
rect 2789 20961 2823 20995
rect 5641 20961 5675 20995
rect 7757 20961 7791 20995
rect 8217 20961 8251 20995
rect 9413 20961 9447 20995
rect 9505 20961 9539 20995
rect 19625 20961 19659 20995
rect 1409 20893 1443 20927
rect 1869 20893 1903 20927
rect 2421 20893 2455 20927
rect 3433 20893 3467 20927
rect 3985 20893 4019 20927
rect 4077 20893 4111 20927
rect 4353 20893 4387 20927
rect 4445 20893 4479 20927
rect 5181 20893 5215 20927
rect 5365 20893 5399 20927
rect 7481 20893 7515 20927
rect 8125 20893 8159 20927
rect 9321 20893 9355 20927
rect 13001 20893 13035 20927
rect 14289 20893 14323 20927
rect 17509 20893 17543 20927
rect 17693 20893 17727 20927
rect 21465 20893 21499 20927
rect 23305 20893 23339 20927
rect 23857 20893 23891 20927
rect 24501 20893 24535 20927
rect 3341 20825 3375 20859
rect 4905 20825 4939 20859
rect 5917 20825 5951 20859
rect 10425 20825 10459 20859
rect 16221 20825 16255 20859
rect 16437 20825 16471 20859
rect 19901 20825 19935 20859
rect 21557 20825 21591 20859
rect 25053 20825 25087 20859
rect 1593 20757 1627 20791
rect 4261 20757 4295 20791
rect 5549 20757 5583 20791
rect 16589 20757 16623 20791
rect 23397 20757 23431 20791
rect 23949 20757 23983 20791
rect 3433 20553 3467 20587
rect 3985 20553 4019 20587
rect 7481 20553 7515 20587
rect 13185 20553 13219 20587
rect 19717 20553 19751 20587
rect 5181 20485 5215 20519
rect 5381 20485 5415 20519
rect 10609 20485 10643 20519
rect 17049 20485 17083 20519
rect 24777 20485 24811 20519
rect 2789 20417 2823 20451
rect 3157 20417 3191 20451
rect 3249 20417 3283 20451
rect 3617 20417 3651 20451
rect 4629 20417 4663 20451
rect 5917 20417 5951 20451
rect 6561 20417 6595 20451
rect 7113 20417 7147 20451
rect 7297 20417 7331 20451
rect 8217 20417 8251 20451
rect 10517 20417 10551 20451
rect 13001 20417 13035 20451
rect 13461 20417 13495 20451
rect 13645 20417 13679 20451
rect 15209 20417 15243 20451
rect 15761 20417 15795 20451
rect 16865 20417 16899 20451
rect 17141 20417 17175 20451
rect 17877 20417 17911 20451
rect 17969 20417 18003 20451
rect 18245 20417 18279 20451
rect 20545 20417 20579 20451
rect 21005 20417 21039 20451
rect 22937 20417 22971 20451
rect 23305 20417 23339 20451
rect 3709 20349 3743 20383
rect 4721 20349 4755 20383
rect 5733 20349 5767 20383
rect 6745 20349 6779 20383
rect 8493 20349 8527 20383
rect 10701 20349 10735 20383
rect 13829 20349 13863 20383
rect 18153 20349 18187 20383
rect 20637 20349 20671 20383
rect 21281 20349 21315 20383
rect 5549 20281 5583 20315
rect 10149 20281 10183 20315
rect 15577 20281 15611 20315
rect 2881 20213 2915 20247
rect 3617 20213 3651 20247
rect 4629 20213 4663 20247
rect 4997 20213 5031 20247
rect 5365 20213 5399 20247
rect 6101 20213 6135 20247
rect 9965 20213 9999 20247
rect 15669 20213 15703 20247
rect 16037 20213 16071 20247
rect 16221 20213 16255 20247
rect 16681 20213 16715 20247
rect 18061 20213 18095 20247
rect 20821 20213 20855 20247
rect 21281 20213 21315 20247
rect 21557 20213 21591 20247
rect 2973 20009 3007 20043
rect 4629 20009 4663 20043
rect 4997 20009 5031 20043
rect 5733 20009 5767 20043
rect 5917 20009 5951 20043
rect 7021 20009 7055 20043
rect 9229 20009 9263 20043
rect 11437 20009 11471 20043
rect 12725 20009 12759 20043
rect 20085 20009 20119 20043
rect 6745 19941 6779 19975
rect 7481 19941 7515 19975
rect 3617 19873 3651 19907
rect 4445 19873 4479 19907
rect 5181 19873 5215 19907
rect 8585 19873 8619 19907
rect 9689 19873 9723 19907
rect 19441 19873 19475 19907
rect 20453 19873 20487 19907
rect 21741 19873 21775 19907
rect 22017 19873 22051 19907
rect 24041 19873 24075 19907
rect 2421 19805 2455 19839
rect 2605 19805 2639 19839
rect 2789 19805 2823 19839
rect 2973 19805 3007 19839
rect 3341 19805 3375 19839
rect 3433 19805 3467 19839
rect 3801 19805 3835 19839
rect 4537 19805 4571 19839
rect 4905 19805 4939 19839
rect 5641 19805 5675 19839
rect 5825 19805 5859 19839
rect 6101 19805 6135 19839
rect 6193 19805 6227 19839
rect 6561 19805 6595 19839
rect 6929 19805 6963 19839
rect 7297 19805 7331 19839
rect 8493 19805 8527 19839
rect 9137 19805 9171 19839
rect 9597 19805 9631 19839
rect 12541 19805 12575 19839
rect 12817 19805 12851 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 16037 19805 16071 19839
rect 16313 19805 16347 19839
rect 16497 19805 16531 19839
rect 16589 19805 16623 19839
rect 16681 19805 16715 19839
rect 17877 19805 17911 19839
rect 18061 19805 18095 19839
rect 19257 19805 19291 19839
rect 20269 19805 20303 19839
rect 20361 19805 20395 19839
rect 20545 19805 20579 19839
rect 20821 19805 20855 19839
rect 21281 19805 21315 19839
rect 21373 19805 21407 19839
rect 3617 19737 3651 19771
rect 8401 19737 8435 19771
rect 9965 19737 9999 19771
rect 16221 19737 16255 19771
rect 21465 19737 21499 19771
rect 21583 19737 21617 19771
rect 22293 19737 22327 19771
rect 2513 19669 2547 19703
rect 3157 19669 3191 19703
rect 5457 19669 5491 19703
rect 6377 19669 6411 19703
rect 8033 19669 8067 19703
rect 9413 19669 9447 19703
rect 12909 19669 12943 19703
rect 14197 19669 14231 19703
rect 15853 19669 15887 19703
rect 16865 19669 16899 19703
rect 18245 19669 18279 19703
rect 20913 19669 20947 19703
rect 21097 19669 21131 19703
rect 3157 19465 3191 19499
rect 4813 19465 4847 19499
rect 8401 19465 8435 19499
rect 13553 19465 13587 19499
rect 13845 19465 13879 19499
rect 14013 19465 14047 19499
rect 16405 19465 16439 19499
rect 17049 19465 17083 19499
rect 18153 19465 18187 19499
rect 20269 19465 20303 19499
rect 20361 19465 20395 19499
rect 22201 19465 22235 19499
rect 23213 19465 23247 19499
rect 1685 19397 1719 19431
rect 11621 19397 11655 19431
rect 13645 19397 13679 19431
rect 17877 19397 17911 19431
rect 18889 19397 18923 19431
rect 19901 19397 19935 19431
rect 20117 19397 20151 19431
rect 22385 19397 22419 19431
rect 1409 19329 1443 19363
rect 3249 19329 3283 19363
rect 3801 19329 3835 19363
rect 3985 19329 4019 19363
rect 4261 19329 4295 19363
rect 6377 19329 6411 19363
rect 6561 19329 6595 19363
rect 8585 19329 8619 19363
rect 9505 19329 9539 19363
rect 9597 19329 9631 19363
rect 11529 19329 11563 19363
rect 11805 19329 11839 19363
rect 15853 19329 15887 19363
rect 16221 19329 16255 19363
rect 17509 19329 17543 19363
rect 17601 19329 17635 19363
rect 18061 19329 18095 19363
rect 18245 19329 18279 19363
rect 18337 19329 18371 19363
rect 19073 19329 19107 19363
rect 20535 19329 20569 19363
rect 20821 19329 20855 19363
rect 21189 19329 21223 19363
rect 21465 19329 21499 19363
rect 21833 19329 21867 19363
rect 22017 19329 22051 19363
rect 22293 19329 22327 19363
rect 23121 19329 23155 19363
rect 3341 19261 3375 19295
rect 4537 19261 4571 19295
rect 9873 19261 9907 19295
rect 12081 19261 12115 19295
rect 15761 19261 15795 19295
rect 17969 19261 18003 19295
rect 18521 19261 18555 19295
rect 20729 19261 20763 19295
rect 21373 19261 21407 19295
rect 4169 19193 4203 19227
rect 9321 19193 9355 19227
rect 16681 19193 16715 19227
rect 17325 19193 17359 19227
rect 20637 19193 20671 19227
rect 21281 19193 21315 19227
rect 3433 19125 3467 19159
rect 3617 19125 3651 19159
rect 3985 19125 4019 19159
rect 4629 19125 4663 19159
rect 6469 19125 6503 19159
rect 11345 19125 11379 19159
rect 13829 19125 13863 19159
rect 16221 19125 16255 19159
rect 17049 19125 17083 19159
rect 17233 19125 17267 19159
rect 19257 19125 19291 19159
rect 20085 19125 20119 19159
rect 21005 19125 21039 19159
rect 2421 18921 2455 18955
rect 6561 18921 6595 18955
rect 7205 18921 7239 18955
rect 9781 18921 9815 18955
rect 10977 18921 11011 18955
rect 14289 18921 14323 18955
rect 19579 18921 19613 18955
rect 20269 18921 20303 18955
rect 20453 18921 20487 18955
rect 23857 18921 23891 18955
rect 14473 18853 14507 18887
rect 16405 18853 16439 18887
rect 7389 18785 7423 18819
rect 10333 18785 10367 18819
rect 13185 18785 13219 18819
rect 15761 18785 15795 18819
rect 20085 18785 20119 18819
rect 21097 18785 21131 18819
rect 2329 18717 2363 18751
rect 4997 18717 5031 18751
rect 7113 18717 7147 18751
rect 10885 18717 10919 18751
rect 12633 18717 12667 18751
rect 13277 18717 13311 18751
rect 14565 18717 14599 18751
rect 15945 18717 15979 18751
rect 16221 18717 16255 18751
rect 17233 18717 17267 18751
rect 17509 18717 17543 18751
rect 17601 18717 17635 18751
rect 17877 18717 17911 18751
rect 18337 18717 18371 18751
rect 18521 18717 18555 18751
rect 19441 18717 19475 18751
rect 19717 18717 19751 18751
rect 19901 18717 19935 18751
rect 20269 18717 20303 18751
rect 20821 18717 20855 18751
rect 20913 18717 20947 18751
rect 21005 18717 21039 18751
rect 21281 18717 21315 18751
rect 21649 18717 21683 18751
rect 22109 18717 22143 18751
rect 23949 18717 23983 18751
rect 5273 18649 5307 18683
rect 10241 18649 10275 18683
rect 13553 18649 13587 18683
rect 14105 18649 14139 18683
rect 14657 18649 14691 18683
rect 16405 18649 16439 18683
rect 17141 18649 17175 18683
rect 17417 18649 17451 18683
rect 18061 18649 18095 18683
rect 19993 18649 20027 18683
rect 21465 18649 21499 18683
rect 21557 18649 21591 18683
rect 22385 18649 22419 18683
rect 24041 18649 24075 18683
rect 5089 18581 5123 18615
rect 7665 18581 7699 18615
rect 10149 18581 10183 18615
rect 14305 18581 14339 18615
rect 16129 18581 16163 18615
rect 16865 18581 16899 18615
rect 16957 18581 16991 18615
rect 17785 18581 17819 18615
rect 18245 18581 18279 18615
rect 18705 18581 18739 18615
rect 19901 18581 19935 18615
rect 20637 18581 20671 18615
rect 21833 18581 21867 18615
rect 2605 18377 2639 18411
rect 2973 18377 3007 18411
rect 4261 18377 4295 18411
rect 7665 18377 7699 18411
rect 8585 18377 8619 18411
rect 14105 18377 14139 18411
rect 16681 18377 16715 18411
rect 17601 18377 17635 18411
rect 17995 18377 18029 18411
rect 20009 18377 20043 18411
rect 20177 18377 20211 18411
rect 20637 18377 20671 18411
rect 21373 18377 21407 18411
rect 25145 18377 25179 18411
rect 6377 18309 6411 18343
rect 8677 18309 8711 18343
rect 10701 18309 10735 18343
rect 16129 18309 16163 18343
rect 16345 18309 16379 18343
rect 17785 18309 17819 18343
rect 19809 18309 19843 18343
rect 2329 18241 2363 18275
rect 3801 18241 3835 18275
rect 4353 18241 4387 18275
rect 4721 18241 4755 18275
rect 5365 18241 5399 18275
rect 5825 18241 5859 18275
rect 6009 18241 6043 18275
rect 6193 18241 6227 18275
rect 9229 18241 9263 18275
rect 10609 18241 10643 18275
rect 10793 18241 10827 18275
rect 10885 18241 10919 18275
rect 11069 18241 11103 18275
rect 11713 18241 11747 18275
rect 11897 18241 11931 18275
rect 12357 18241 12391 18275
rect 12909 18241 12943 18275
rect 13553 18241 13587 18275
rect 13645 18241 13679 18275
rect 13921 18241 13955 18275
rect 14381 18241 14415 18275
rect 14657 18241 14691 18275
rect 14841 18241 14875 18275
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 17417 18241 17451 18275
rect 17693 18241 17727 18275
rect 20821 18241 20855 18275
rect 21005 18241 21039 18275
rect 21097 18241 21131 18275
rect 21189 18241 21223 18275
rect 21373 18241 21407 18275
rect 25053 18241 25087 18275
rect 3065 18173 3099 18207
rect 3249 18173 3283 18207
rect 4445 18173 4479 18207
rect 4997 18173 5031 18207
rect 5457 18173 5491 18207
rect 8769 18173 8803 18207
rect 11253 18173 11287 18207
rect 11529 18173 11563 18207
rect 11805 18173 11839 18207
rect 11989 18173 12023 18207
rect 12173 18173 12207 18207
rect 14197 18173 14231 18207
rect 17141 18173 17175 18207
rect 3893 18105 3927 18139
rect 5273 18105 5307 18139
rect 8217 18105 8251 18139
rect 11161 18105 11195 18139
rect 12541 18105 12575 18139
rect 16497 18105 16531 18139
rect 18153 18105 18187 18139
rect 2145 18037 2179 18071
rect 3617 18037 3651 18071
rect 4813 18037 4847 18071
rect 5365 18037 5399 18071
rect 5733 18037 5767 18071
rect 9045 18037 9079 18071
rect 11253 18037 11287 18071
rect 13185 18037 13219 18071
rect 13369 18037 13403 18071
rect 13829 18037 13863 18071
rect 14565 18037 14599 18071
rect 14749 18037 14783 18071
rect 16313 18037 16347 18071
rect 17049 18037 17083 18071
rect 17969 18037 18003 18071
rect 19993 18037 20027 18071
rect 6101 17833 6135 17867
rect 6929 17833 6963 17867
rect 13093 17833 13127 17867
rect 13277 17833 13311 17867
rect 13737 17833 13771 17867
rect 14289 17833 14323 17867
rect 16865 17833 16899 17867
rect 7389 17765 7423 17799
rect 7573 17765 7607 17799
rect 12541 17765 12575 17799
rect 3801 17697 3835 17731
rect 6745 17697 6779 17731
rect 8125 17697 8159 17731
rect 12081 17697 12115 17731
rect 19533 17697 19567 17731
rect 23489 17697 23523 17731
rect 1409 17629 1443 17663
rect 3433 17629 3467 17663
rect 5733 17629 5767 17663
rect 6837 17629 6871 17663
rect 7113 17629 7147 17663
rect 8585 17629 8619 17663
rect 8953 17629 8987 17663
rect 9965 17629 9999 17663
rect 10425 17629 10459 17663
rect 14565 17629 14599 17663
rect 17049 17629 17083 17663
rect 17233 17629 17267 17663
rect 17325 17629 17359 17663
rect 17509 17629 17543 17663
rect 19717 17629 19751 17663
rect 21097 17629 21131 17663
rect 21465 17629 21499 17663
rect 22661 17629 22695 17663
rect 23213 17629 23247 17663
rect 1685 17561 1719 17595
rect 4077 17561 4111 17595
rect 6377 17561 6411 17595
rect 6561 17561 6595 17595
rect 8401 17561 8435 17595
rect 10149 17561 10183 17595
rect 12265 17561 12299 17595
rect 12909 17561 12943 17595
rect 13369 17561 13403 17595
rect 13553 17561 13587 17595
rect 14105 17561 14139 17595
rect 18153 17561 18187 17595
rect 20637 17561 20671 17595
rect 20821 17561 20855 17595
rect 21005 17561 21039 17595
rect 21281 17561 21315 17595
rect 21373 17561 21407 17595
rect 5549 17493 5583 17527
rect 6101 17493 6135 17527
rect 6285 17493 6319 17527
rect 7941 17493 7975 17527
rect 8033 17493 8067 17527
rect 8769 17493 8803 17527
rect 9045 17493 9079 17527
rect 10333 17493 10367 17527
rect 12725 17493 12759 17527
rect 13109 17493 13143 17527
rect 14305 17493 14339 17527
rect 14473 17493 14507 17527
rect 14749 17493 14783 17527
rect 19901 17493 19935 17527
rect 21649 17493 21683 17527
rect 22753 17493 22787 17527
rect 2513 17289 2547 17323
rect 9321 17289 9355 17323
rect 10425 17289 10459 17323
rect 11529 17289 11563 17323
rect 18429 17289 18463 17323
rect 21557 17289 21591 17323
rect 2237 17221 2271 17255
rect 6377 17221 6411 17255
rect 6577 17221 6611 17255
rect 13921 17221 13955 17255
rect 14121 17221 14155 17255
rect 16405 17221 16439 17255
rect 16957 17221 16991 17255
rect 22293 17221 22327 17255
rect 24041 17221 24075 17255
rect 2145 17153 2179 17187
rect 2421 17153 2455 17187
rect 4445 17153 4479 17187
rect 6837 17153 6871 17187
rect 7573 17153 7607 17187
rect 10609 17153 10643 17187
rect 10701 17153 10735 17187
rect 10885 17153 10919 17187
rect 10977 17153 11011 17187
rect 11713 17153 11747 17187
rect 14565 17153 14599 17187
rect 14841 17153 14875 17187
rect 16313 17153 16347 17187
rect 19625 17153 19659 17187
rect 20453 17153 20487 17187
rect 22017 17153 22051 17187
rect 25697 17153 25731 17187
rect 4721 17085 4755 17119
rect 6193 17085 6227 17119
rect 7113 17085 7147 17119
rect 7849 17085 7883 17119
rect 9873 17085 9907 17119
rect 11805 17085 11839 17119
rect 11897 17085 11931 17119
rect 11989 17085 12023 17119
rect 16681 17085 16715 17119
rect 19717 17085 19751 17119
rect 19993 17085 20027 17119
rect 20545 17085 20579 17119
rect 20821 17085 20855 17119
rect 21005 17085 21039 17119
rect 10149 17017 10183 17051
rect 14289 17017 14323 17051
rect 25881 17017 25915 17051
rect 6561 16949 6595 16983
rect 6745 16949 6779 16983
rect 6929 16949 6963 16983
rect 7389 16949 7423 16983
rect 10333 16949 10367 16983
rect 14105 16949 14139 16983
rect 14749 16949 14783 16983
rect 15025 16949 15059 16983
rect 1409 16745 1443 16779
rect 4629 16745 4663 16779
rect 4997 16745 5031 16779
rect 8769 16745 8803 16779
rect 13921 16745 13955 16779
rect 10701 16677 10735 16711
rect 19809 16677 19843 16711
rect 23213 16677 23247 16711
rect 4629 16609 4663 16643
rect 5917 16609 5951 16643
rect 7021 16609 7055 16643
rect 11161 16609 11195 16643
rect 11437 16609 11471 16643
rect 12173 16609 12207 16643
rect 20177 16609 20211 16643
rect 21465 16609 21499 16643
rect 1593 16541 1627 16575
rect 4353 16541 4387 16575
rect 5181 16541 5215 16575
rect 5641 16541 5675 16575
rect 6101 16541 6135 16575
rect 6193 16541 6227 16575
rect 8953 16541 8987 16575
rect 9781 16541 9815 16575
rect 9873 16541 9907 16575
rect 10057 16541 10091 16575
rect 10205 16541 10239 16575
rect 10522 16541 10556 16575
rect 11529 16541 11563 16575
rect 11897 16541 11931 16575
rect 12081 16541 12115 16575
rect 14105 16541 14139 16575
rect 17233 16541 17267 16575
rect 17325 16541 17359 16575
rect 19809 16541 19843 16575
rect 19993 16541 20027 16575
rect 20085 16541 20119 16575
rect 20269 16541 20303 16575
rect 20545 16541 20579 16575
rect 20729 16541 20763 16575
rect 21189 16541 21223 16575
rect 21281 16541 21315 16575
rect 23397 16541 23431 16575
rect 7297 16473 7331 16507
rect 9045 16473 9079 16507
rect 10333 16473 10367 16507
rect 10425 16473 10459 16507
rect 12449 16473 12483 16507
rect 14197 16473 14231 16507
rect 20361 16473 20395 16507
rect 21005 16473 21039 16507
rect 21741 16473 21775 16507
rect 4905 16405 4939 16439
rect 5273 16405 5307 16439
rect 5733 16405 5767 16439
rect 21103 16405 21137 16439
rect 23489 16405 23523 16439
rect 3341 16201 3375 16235
rect 3709 16201 3743 16235
rect 5365 16201 5399 16235
rect 6837 16201 6871 16235
rect 8217 16201 8251 16235
rect 10517 16201 10551 16235
rect 12725 16201 12759 16235
rect 13461 16201 13495 16235
rect 20361 16201 20395 16235
rect 21557 16201 21591 16235
rect 12357 16133 12391 16167
rect 12449 16133 12483 16167
rect 19073 16133 19107 16167
rect 21833 16133 21867 16167
rect 2329 16065 2363 16099
rect 2421 16065 2455 16099
rect 2881 16065 2915 16099
rect 2973 16065 3007 16099
rect 6745 16065 6779 16099
rect 8125 16065 8159 16099
rect 8401 16065 8435 16099
rect 10241 16065 10275 16099
rect 10333 16065 10367 16099
rect 12173 16065 12207 16099
rect 12541 16065 12575 16099
rect 13277 16065 13311 16099
rect 16957 16065 16991 16099
rect 22017 16065 22051 16099
rect 22109 16065 22143 16099
rect 3801 15997 3835 16031
rect 3985 15997 4019 16031
rect 5457 15997 5491 16031
rect 5549 15997 5583 16031
rect 6929 15997 6963 16031
rect 7573 15997 7607 16031
rect 10517 15997 10551 16031
rect 13093 15997 13127 16031
rect 17233 15997 17267 16031
rect 18981 15997 19015 16031
rect 21005 15997 21039 16031
rect 2513 15929 2547 15963
rect 21833 15929 21867 15963
rect 2145 15861 2179 15895
rect 2697 15861 2731 15895
rect 3065 15861 3099 15895
rect 4997 15861 5031 15895
rect 6377 15861 6411 15895
rect 3801 15657 3835 15691
rect 11897 15657 11931 15691
rect 16497 15657 16531 15691
rect 17785 15657 17819 15691
rect 18153 15657 18187 15691
rect 22155 15657 22189 15691
rect 3341 15589 3375 15623
rect 1593 15521 1627 15555
rect 1869 15521 1903 15555
rect 4445 15521 4479 15555
rect 7665 15521 7699 15555
rect 16037 15521 16071 15555
rect 16865 15521 16899 15555
rect 17141 15521 17175 15555
rect 19441 15521 19475 15555
rect 20361 15521 20395 15555
rect 4169 15453 4203 15487
rect 5273 15453 5307 15487
rect 7573 15453 7607 15487
rect 7941 15453 7975 15487
rect 8953 15453 8987 15487
rect 9873 15453 9907 15487
rect 10057 15453 10091 15487
rect 10333 15453 10367 15487
rect 12081 15453 12115 15487
rect 13553 15453 13587 15487
rect 15577 15453 15611 15487
rect 16129 15453 16163 15487
rect 16773 15453 16807 15487
rect 17233 15453 17267 15487
rect 17601 15453 17635 15487
rect 18061 15453 18095 15487
rect 19257 15453 19291 15487
rect 20729 15453 20763 15487
rect 7481 15385 7515 15419
rect 17417 15385 17451 15419
rect 17509 15385 17543 15419
rect 4261 15317 4295 15351
rect 6561 15317 6595 15351
rect 7113 15317 7147 15351
rect 8033 15317 8067 15351
rect 9597 15317 9631 15351
rect 9689 15317 9723 15351
rect 10149 15317 10183 15351
rect 10425 15317 10459 15351
rect 13737 15317 13771 15351
rect 15669 15317 15703 15351
rect 8125 15113 8159 15147
rect 11897 15113 11931 15147
rect 11989 15113 12023 15147
rect 13921 15113 13955 15147
rect 17049 15113 17083 15147
rect 20821 15113 20855 15147
rect 1685 15045 1719 15079
rect 8769 15045 8803 15079
rect 9505 15045 9539 15079
rect 12633 15045 12667 15079
rect 16681 15045 16715 15079
rect 1409 14977 1443 15011
rect 4169 14977 4203 15011
rect 6377 14977 6411 15011
rect 11713 14977 11747 15011
rect 12173 14977 12207 15011
rect 12541 14977 12575 15011
rect 16865 14977 16899 15011
rect 17785 14977 17819 15011
rect 18061 14977 18095 15011
rect 18705 14977 18739 15011
rect 18889 14977 18923 15011
rect 19993 14977 20027 15011
rect 20269 14977 20303 15011
rect 20729 14977 20763 15011
rect 4445 14909 4479 14943
rect 6193 14909 6227 14943
rect 6653 14909 6687 14943
rect 8861 14909 8895 14943
rect 8953 14909 8987 14943
rect 9229 14909 9263 14943
rect 11529 14909 11563 14943
rect 14473 14909 14507 14943
rect 14749 14909 14783 14943
rect 16221 14909 16255 14943
rect 17877 14841 17911 14875
rect 3157 14773 3191 14807
rect 8401 14773 8435 14807
rect 10977 14773 11011 14807
rect 12357 14773 12391 14807
rect 18153 14773 18187 14807
rect 19073 14773 19107 14807
rect 20085 14773 20119 14807
rect 20361 14773 20395 14807
rect 4905 14569 4939 14603
rect 5733 14569 5767 14603
rect 6377 14569 6411 14603
rect 6837 14569 6871 14603
rect 11713 14569 11747 14603
rect 13921 14569 13955 14603
rect 14473 14569 14507 14603
rect 17233 14569 17267 14603
rect 8769 14501 8803 14535
rect 11069 14501 11103 14535
rect 16221 14501 16255 14535
rect 7021 14433 7055 14467
rect 9229 14433 9263 14467
rect 10977 14433 11011 14467
rect 12173 14433 12207 14467
rect 12449 14433 12483 14467
rect 14657 14433 14691 14467
rect 16681 14433 16715 14467
rect 18245 14433 18279 14467
rect 19257 14433 19291 14467
rect 4261 14365 4295 14399
rect 5089 14365 5123 14399
rect 5641 14365 5675 14399
rect 6561 14365 6595 14399
rect 6745 14365 6779 14399
rect 9137 14365 9171 14399
rect 11253 14365 11287 14399
rect 11345 14365 11379 14399
rect 11529 14365 11563 14399
rect 14565 14365 14599 14399
rect 15117 14365 15151 14399
rect 15393 14365 15427 14399
rect 16129 14365 16163 14399
rect 16497 14365 16531 14399
rect 17325 14365 17359 14399
rect 17509 14365 17543 14399
rect 17693 14365 17727 14399
rect 18521 14365 18555 14399
rect 18705 14365 18739 14399
rect 18823 14365 18857 14399
rect 18981 14365 19015 14399
rect 7297 14297 7331 14331
rect 9505 14297 9539 14331
rect 14105 14297 14139 14331
rect 14289 14297 14323 14331
rect 15761 14297 15795 14331
rect 15945 14297 15979 14331
rect 16221 14297 16255 14331
rect 17417 14297 17451 14331
rect 18613 14297 18647 14331
rect 19533 14297 19567 14331
rect 21281 14297 21315 14331
rect 4813 14229 4847 14263
rect 8953 14229 8987 14263
rect 15215 14229 15249 14263
rect 15301 14229 15335 14263
rect 16405 14229 16439 14263
rect 18337 14229 18371 14263
rect 6653 14025 6687 14059
rect 7389 14025 7423 14059
rect 8493 14025 8527 14059
rect 11161 14025 11195 14059
rect 13645 14025 13679 14059
rect 17969 14025 18003 14059
rect 18613 14025 18647 14059
rect 5089 13957 5123 13991
rect 5273 13957 5307 13991
rect 8861 13957 8895 13991
rect 8953 13957 8987 13991
rect 12173 13957 12207 13991
rect 13829 13957 13863 13991
rect 17049 13957 17083 13991
rect 17249 13957 17283 13991
rect 17601 13957 17635 13991
rect 17817 13957 17851 13991
rect 4445 13889 4479 13923
rect 4721 13889 4755 13923
rect 5733 13889 5767 13923
rect 5917 13889 5951 13923
rect 6469 13889 6503 13923
rect 7021 13889 7055 13923
rect 7113 13889 7147 13923
rect 7573 13889 7607 13923
rect 9321 13889 9355 13923
rect 10977 13889 11011 13923
rect 13737 13889 13771 13923
rect 18245 13889 18279 13923
rect 18889 13889 18923 13923
rect 6101 13821 6135 13855
rect 9045 13821 9079 13855
rect 9597 13821 9631 13855
rect 10793 13821 10827 13855
rect 11897 13821 11931 13855
rect 18153 13821 18187 13855
rect 19257 13821 19291 13855
rect 4261 13753 4295 13787
rect 17417 13753 17451 13787
rect 4629 13685 4663 13719
rect 6009 13685 6043 13719
rect 6101 13685 6135 13719
rect 7297 13685 7331 13719
rect 17233 13685 17267 13719
rect 17785 13685 17819 13719
rect 20683 13685 20717 13719
rect 6561 13481 6595 13515
rect 6745 13481 6779 13515
rect 7113 13481 7147 13515
rect 7573 13481 7607 13515
rect 12541 13481 12575 13515
rect 16405 13481 16439 13515
rect 17877 13481 17911 13515
rect 19901 13481 19935 13515
rect 20361 13481 20395 13515
rect 25973 13481 26007 13515
rect 5181 13413 5215 13447
rect 6009 13413 6043 13447
rect 7757 13413 7791 13447
rect 16313 13413 16347 13447
rect 18153 13413 18187 13447
rect 20545 13413 20579 13447
rect 5365 13345 5399 13379
rect 11345 13345 11379 13379
rect 15853 13345 15887 13379
rect 17325 13345 17359 13379
rect 18245 13345 18279 13379
rect 18521 13345 18555 13379
rect 19257 13345 19291 13379
rect 20821 13345 20855 13379
rect 3801 13277 3835 13311
rect 6285 13277 6319 13311
rect 6377 13277 6411 13311
rect 6653 13277 6687 13311
rect 10609 13277 10643 13311
rect 12173 13277 12207 13311
rect 12357 13277 12391 13311
rect 12817 13277 12851 13311
rect 14105 13277 14139 13311
rect 16037 13277 16071 13311
rect 16129 13277 16163 13311
rect 16405 13277 16439 13311
rect 16589 13277 16623 13311
rect 16681 13277 16715 13311
rect 16865 13277 16899 13311
rect 17049 13277 17083 13311
rect 17509 13277 17543 13311
rect 17785 13277 17819 13311
rect 18061 13277 18095 13311
rect 18337 13277 18371 13311
rect 18705 13277 18739 13311
rect 18797 13277 18831 13311
rect 18889 13277 18923 13311
rect 18981 13277 19015 13311
rect 19993 13277 20027 13311
rect 20269 13277 20303 13311
rect 25789 13277 25823 13311
rect 4068 13209 4102 13243
rect 5917 13209 5951 13243
rect 7389 13209 7423 13243
rect 10793 13209 10827 13243
rect 10977 13209 11011 13243
rect 14381 13209 14415 13243
rect 16957 13209 16991 13243
rect 17693 13209 17727 13243
rect 21097 13209 21131 13243
rect 6193 13141 6227 13175
rect 7589 13141 7623 13175
rect 11897 13141 11931 13175
rect 12909 13141 12943 13175
rect 17233 13141 17267 13175
rect 22569 13141 22603 13175
rect 3525 12937 3559 12971
rect 5181 12937 5215 12971
rect 13599 12937 13633 12971
rect 15393 12937 15427 12971
rect 16681 12937 16715 12971
rect 18613 12937 18647 12971
rect 21097 12937 21131 12971
rect 23121 12937 23155 12971
rect 1501 12869 1535 12903
rect 10885 12869 10919 12903
rect 2401 12801 2435 12835
rect 3801 12801 3835 12835
rect 4068 12801 4102 12835
rect 5273 12801 5307 12835
rect 7113 12801 7147 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 8033 12801 8067 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10149 12801 10183 12835
rect 10609 12801 10643 12835
rect 11069 12801 11103 12835
rect 11529 12801 11563 12835
rect 11805 12801 11839 12835
rect 15301 12801 15335 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 17601 12801 17635 12835
rect 18797 12801 18831 12835
rect 19073 12801 19107 12835
rect 21373 12801 21407 12835
rect 21465 12801 21499 12835
rect 22661 12801 22695 12835
rect 22753 12801 22787 12835
rect 23029 12801 23063 12835
rect 2145 12733 2179 12767
rect 6469 12733 6503 12767
rect 8125 12733 8159 12767
rect 10333 12733 10367 12767
rect 10425 12733 10459 12767
rect 11253 12733 11287 12767
rect 12173 12733 12207 12767
rect 16865 12733 16899 12767
rect 16957 12733 16991 12767
rect 17141 12733 17175 12767
rect 17509 12733 17543 12767
rect 21281 12733 21315 12767
rect 21557 12733 21591 12767
rect 22017 12733 22051 12767
rect 9597 12665 9631 12699
rect 10241 12665 10275 12699
rect 18889 12665 18923 12699
rect 18981 12665 19015 12699
rect 1593 12597 1627 12631
rect 5917 12597 5951 12631
rect 7021 12597 7055 12631
rect 7113 12597 7147 12631
rect 8769 12597 8803 12631
rect 10793 12597 10827 12631
rect 11713 12597 11747 12631
rect 17325 12597 17359 12631
rect 17785 12597 17819 12631
rect 22845 12597 22879 12631
rect 3525 12393 3559 12427
rect 6561 12393 6595 12427
rect 10977 12393 11011 12427
rect 13599 12393 13633 12427
rect 16681 12393 16715 12427
rect 17141 12393 17175 12427
rect 4813 12325 4847 12359
rect 8493 12325 8527 12359
rect 16543 12325 16577 12359
rect 1777 12257 1811 12291
rect 2145 12257 2179 12291
rect 3801 12257 3835 12291
rect 7021 12257 7055 12291
rect 10425 12257 10459 12291
rect 11713 12257 11747 12291
rect 12173 12257 12207 12291
rect 16313 12257 16347 12291
rect 16773 12257 16807 12291
rect 1685 12189 1719 12223
rect 4721 12189 4755 12223
rect 5089 12189 5123 12223
rect 5917 12189 5951 12223
rect 6065 12189 6099 12223
rect 6285 12189 6319 12223
rect 6382 12189 6416 12223
rect 6653 12189 6687 12223
rect 7288 12189 7322 12223
rect 8493 12189 8527 12223
rect 8769 12189 8803 12223
rect 9321 12189 9355 12223
rect 11161 12189 11195 12223
rect 11805 12189 11839 12223
rect 15025 12189 15059 12223
rect 15761 12189 15795 12223
rect 16405 12189 16439 12223
rect 16865 12189 16899 12223
rect 17049 12189 17083 12223
rect 17233 12189 17267 12223
rect 20729 12189 20763 12223
rect 24409 12189 24443 12223
rect 2412 12121 2446 12155
rect 6193 12121 6227 12155
rect 8677 12121 8711 12155
rect 21005 12121 21039 12155
rect 22753 12121 22787 12155
rect 2053 12053 2087 12087
rect 4445 12053 4479 12087
rect 5641 12053 5675 12087
rect 6837 12053 6871 12087
rect 8401 12053 8435 12087
rect 9965 12053 9999 12087
rect 15117 12053 15151 12087
rect 24501 12053 24535 12087
rect 2329 11849 2363 11883
rect 2697 11849 2731 11883
rect 4353 11849 4387 11883
rect 5825 11849 5859 11883
rect 6377 11849 6411 11883
rect 7205 11849 7239 11883
rect 8309 11849 8343 11883
rect 9137 11849 9171 11883
rect 11023 11849 11057 11883
rect 11897 11849 11931 11883
rect 13185 11849 13219 11883
rect 18813 11849 18847 11883
rect 20913 11849 20947 11883
rect 21833 11849 21867 11883
rect 2145 11781 2179 11815
rect 2513 11781 2547 11815
rect 2973 11781 3007 11815
rect 5549 11781 5583 11815
rect 7113 11781 7147 11815
rect 7573 11781 7607 11815
rect 14565 11781 14599 11815
rect 16313 11781 16347 11815
rect 17049 11781 17083 11815
rect 18613 11781 18647 11815
rect 22661 11781 22695 11815
rect 2421 11713 2455 11747
rect 2789 11713 2823 11747
rect 2881 11713 2915 11747
rect 3065 11713 3099 11747
rect 3249 11713 3283 11747
rect 3433 11713 3467 11747
rect 3801 11713 3835 11747
rect 4294 11713 4328 11747
rect 4721 11713 4755 11747
rect 5181 11713 5215 11747
rect 5329 11713 5363 11747
rect 5457 11713 5491 11747
rect 5646 11713 5680 11747
rect 6544 11713 6578 11747
rect 6654 11713 6688 11747
rect 6929 11713 6963 11747
rect 7481 11713 7515 11747
rect 9597 11713 9631 11747
rect 11161 11713 11195 11747
rect 11529 11713 11563 11747
rect 11897 11713 11931 11747
rect 12173 11713 12207 11747
rect 13093 11713 13127 11747
rect 14289 11713 14323 11747
rect 16221 11713 16255 11747
rect 16773 11713 16807 11747
rect 20453 11713 20487 11747
rect 21097 11713 21131 11747
rect 21189 11713 21223 11747
rect 21281 11713 21315 11747
rect 21399 11713 21433 11747
rect 22017 11713 22051 11747
rect 22109 11713 22143 11747
rect 22293 11713 22327 11747
rect 22477 11713 22511 11747
rect 23121 11713 23155 11747
rect 24961 11713 24995 11747
rect 25053 11713 25087 11747
rect 3617 11645 3651 11679
rect 4813 11645 4847 11679
rect 7389 11645 7423 11679
rect 7665 11645 7699 11679
rect 8585 11645 8619 11679
rect 9229 11645 9263 11679
rect 11253 11645 11287 11679
rect 11805 11645 11839 11679
rect 12449 11645 12483 11679
rect 20545 11645 20579 11679
rect 21557 11645 21591 11679
rect 22845 11645 22879 11679
rect 23489 11645 23523 11679
rect 2145 11577 2179 11611
rect 2513 11577 2547 11611
rect 3893 11577 3927 11611
rect 4169 11577 4203 11611
rect 20821 11577 20855 11611
rect 22201 11577 22235 11611
rect 6837 11509 6871 11543
rect 11621 11509 11655 11543
rect 16037 11509 16071 11543
rect 18521 11509 18555 11543
rect 18797 11509 18831 11543
rect 18981 11509 19015 11543
rect 25697 11509 25731 11543
rect 3893 11305 3927 11339
rect 4905 11305 4939 11339
rect 5457 11305 5491 11339
rect 5641 11305 5675 11339
rect 6009 11305 6043 11339
rect 6561 11305 6595 11339
rect 8769 11305 8803 11339
rect 11023 11305 11057 11339
rect 11621 11305 11655 11339
rect 12173 11305 12207 11339
rect 15669 11305 15703 11339
rect 17877 11305 17911 11339
rect 20913 11305 20947 11339
rect 21925 11305 21959 11339
rect 22845 11305 22879 11339
rect 24041 11305 24075 11339
rect 4721 11237 4755 11271
rect 5273 11237 5307 11271
rect 6377 11237 6411 11271
rect 11345 11237 11379 11271
rect 15853 11237 15887 11271
rect 19257 11237 19291 11271
rect 21097 11237 21131 11271
rect 22385 11237 22419 11271
rect 23673 11237 23707 11271
rect 24409 11237 24443 11271
rect 4997 11169 5031 11203
rect 6101 11169 6135 11203
rect 9597 11169 9631 11203
rect 11621 11169 11655 11203
rect 18245 11169 18279 11203
rect 18337 11169 18371 11203
rect 19717 11169 19751 11203
rect 22109 11169 22143 11203
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4445 11101 4479 11135
rect 5549 11101 5583 11135
rect 7389 11101 7423 11135
rect 9229 11101 9263 11135
rect 11253 11101 11287 11135
rect 11529 11101 11563 11135
rect 11897 11101 11931 11135
rect 13737 11101 13771 11135
rect 13921 11101 13955 11135
rect 14197 11101 14231 11135
rect 14565 11101 14599 11135
rect 14841 11101 14875 11135
rect 15025 11101 15059 11135
rect 17785 11101 17819 11135
rect 18429 11101 18463 11135
rect 18521 11101 18555 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 19809 11101 19843 11135
rect 21373 11101 21407 11135
rect 21465 11101 21499 11135
rect 21557 11101 21591 11135
rect 21649 11101 21683 11135
rect 21833 11101 21867 11135
rect 22477 11101 22511 11135
rect 22753 11101 22787 11135
rect 23673 11101 23707 11135
rect 23949 11101 23983 11135
rect 24041 11101 24075 11135
rect 24225 11101 24259 11135
rect 24409 11101 24443 11135
rect 24685 11101 24719 11135
rect 6745 11033 6779 11067
rect 7656 11033 7690 11067
rect 14381 11033 14415 11067
rect 14473 11033 14507 11067
rect 15485 11033 15519 11067
rect 15701 11033 15735 11067
rect 20729 11033 20763 11067
rect 20945 11033 20979 11067
rect 22569 11033 22603 11067
rect 23857 11033 23891 11067
rect 6837 10965 6871 10999
rect 13829 10965 13863 10999
rect 14749 10965 14783 10999
rect 14933 10965 14967 10999
rect 18061 10965 18095 10999
rect 21189 10965 21223 10999
rect 24593 10965 24627 10999
rect 6577 10761 6611 10795
rect 9137 10761 9171 10795
rect 11713 10761 11747 10795
rect 18245 10761 18279 10795
rect 22201 10761 22235 10795
rect 24041 10761 24075 10795
rect 2421 10693 2455 10727
rect 2637 10693 2671 10727
rect 6377 10693 6411 10727
rect 19349 10693 19383 10727
rect 21281 10693 21315 10727
rect 21833 10693 21867 10727
rect 24317 10693 24351 10727
rect 25145 10693 25179 10727
rect 4445 10625 4479 10659
rect 8677 10625 8711 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 11529 10625 11563 10659
rect 13553 10625 13587 10659
rect 13737 10625 13771 10659
rect 13829 10625 13863 10659
rect 15761 10625 15795 10659
rect 18429 10625 18463 10659
rect 18521 10625 18555 10659
rect 18797 10625 18831 10659
rect 18889 10625 18923 10659
rect 19073 10625 19107 10659
rect 19533 10625 19567 10659
rect 19625 10625 19659 10659
rect 21097 10625 21131 10659
rect 21373 10625 21407 10659
rect 21465 10625 21499 10659
rect 22017 10625 22051 10659
rect 22293 10625 22327 10659
rect 23673 10625 23707 10659
rect 23857 10625 23891 10659
rect 24133 10625 24167 10659
rect 24409 10625 24443 10659
rect 24501 10625 24535 10659
rect 24777 10625 24811 10659
rect 24961 10625 24995 10659
rect 5549 10557 5583 10591
rect 8769 10557 8803 10591
rect 6745 10489 6779 10523
rect 19349 10489 19383 10523
rect 2605 10421 2639 10455
rect 2789 10421 2823 10455
rect 4997 10421 5031 10455
rect 6193 10421 6227 10455
rect 6561 10421 6595 10455
rect 13553 10421 13587 10455
rect 13921 10421 13955 10455
rect 15853 10421 15887 10455
rect 18705 10421 18739 10455
rect 19257 10421 19291 10455
rect 21649 10421 21683 10455
rect 24685 10421 24719 10455
rect 7297 10217 7331 10251
rect 9137 10217 9171 10251
rect 11989 10217 12023 10251
rect 14381 10217 14415 10251
rect 15945 10217 15979 10251
rect 16405 10217 16439 10251
rect 17693 10217 17727 10251
rect 18429 10217 18463 10251
rect 19625 10217 19659 10251
rect 20407 10217 20441 10251
rect 22845 10217 22879 10251
rect 23029 10217 23063 10251
rect 24225 10217 24259 10251
rect 24961 10217 24995 10251
rect 16865 10149 16899 10183
rect 17325 10149 17359 10183
rect 17877 10149 17911 10183
rect 20545 10149 20579 10183
rect 25053 10149 25087 10183
rect 2237 10081 2271 10115
rect 20821 10081 20855 10115
rect 21097 10081 21131 10115
rect 23949 10081 23983 10115
rect 24501 10081 24535 10115
rect 2145 10013 2179 10047
rect 4997 10013 5031 10047
rect 5181 10013 5215 10047
rect 5273 10013 5307 10047
rect 7757 10013 7791 10047
rect 9045 10013 9079 10047
rect 9229 10013 9263 10047
rect 11437 10013 11471 10047
rect 12541 10013 12575 10047
rect 12633 10013 12667 10047
rect 12725 10013 12759 10047
rect 12909 10013 12943 10047
rect 13185 10013 13219 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 15117 10013 15151 10047
rect 16681 10013 16715 10047
rect 18429 10013 18463 10047
rect 18521 10013 18555 10047
rect 19257 10013 19291 10047
rect 20269 10013 20303 10047
rect 20729 10013 20763 10047
rect 23305 10013 23339 10047
rect 23397 10013 23431 10047
rect 23857 10013 23891 10047
rect 24593 10013 24627 10047
rect 25053 10013 25087 10047
rect 25237 10013 25271 10047
rect 25329 10013 25363 10047
rect 2482 9945 2516 9979
rect 7113 9945 7147 9979
rect 7313 9945 7347 9979
rect 13369 9945 13403 9979
rect 14105 9945 14139 9979
rect 15301 9945 15335 9979
rect 15761 9945 15795 9979
rect 15977 9945 16011 9979
rect 16313 9945 16347 9979
rect 19441 9945 19475 9979
rect 22661 9945 22695 9979
rect 22877 9945 22911 9979
rect 23581 9945 23615 9979
rect 1961 9877 1995 9911
rect 3617 9877 3651 9911
rect 5181 9877 5215 9911
rect 6561 9877 6595 9911
rect 7481 9877 7515 9911
rect 7573 9877 7607 9911
rect 12265 9877 12299 9911
rect 13737 9877 13771 9911
rect 14565 9877 14599 9911
rect 16129 9877 16163 9911
rect 17693 9877 17727 9911
rect 18797 9877 18831 9911
rect 20729 9877 20763 9911
rect 22569 9877 22603 9911
rect 25421 9877 25455 9911
rect 9689 9673 9723 9707
rect 14105 9673 14139 9707
rect 16773 9673 16807 9707
rect 6009 9605 6043 9639
rect 11989 9605 12023 9639
rect 12449 9605 12483 9639
rect 13553 9605 13587 9639
rect 14473 9605 14507 9639
rect 15301 9605 15335 9639
rect 15761 9605 15795 9639
rect 17141 9605 17175 9639
rect 17341 9605 17375 9639
rect 17601 9605 17635 9639
rect 17801 9605 17835 9639
rect 18429 9605 18463 9639
rect 18705 9605 18739 9639
rect 19441 9605 19475 9639
rect 20729 9605 20763 9639
rect 23857 9605 23891 9639
rect 1777 9537 1811 9571
rect 2237 9537 2271 9571
rect 2493 9537 2527 9571
rect 4077 9537 4111 9571
rect 4629 9537 4663 9571
rect 4777 9537 4811 9571
rect 4905 9537 4939 9571
rect 4997 9537 5031 9571
rect 5135 9537 5169 9571
rect 6377 9537 6411 9571
rect 6644 9537 6678 9571
rect 8033 9537 8067 9571
rect 8309 9537 8343 9571
rect 8565 9537 8599 9571
rect 10149 9537 10183 9571
rect 10241 9537 10275 9571
rect 11897 9537 11931 9571
rect 12357 9537 12391 9571
rect 12541 9537 12575 9571
rect 12909 9537 12943 9571
rect 13277 9537 13311 9571
rect 13737 9537 13771 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 14289 9537 14323 9571
rect 14565 9537 14599 9571
rect 14933 9537 14967 9571
rect 16037 9537 16071 9571
rect 16773 9537 16807 9571
rect 16865 9537 16899 9571
rect 18061 9537 18095 9571
rect 18889 9537 18923 9571
rect 18981 9537 19015 9571
rect 19165 9537 19199 9571
rect 19257 9537 19291 9571
rect 19349 9537 19383 9571
rect 21005 9537 21039 9571
rect 21373 9537 21407 9571
rect 21557 9537 21591 9571
rect 22017 9537 22051 9571
rect 22109 9537 22143 9571
rect 22293 9537 22327 9571
rect 1869 9469 1903 9503
rect 5365 9469 5399 9503
rect 10425 9469 10459 9503
rect 12081 9469 12115 9503
rect 12817 9469 12851 9503
rect 15945 9469 15979 9503
rect 20821 9469 20855 9503
rect 21465 9469 21499 9503
rect 22201 9469 22235 9503
rect 23581 9469 23615 9503
rect 25605 9469 25639 9503
rect 5273 9401 5307 9435
rect 7849 9401 7883 9435
rect 13461 9401 13495 9435
rect 16221 9401 16255 9435
rect 18613 9401 18647 9435
rect 2053 9333 2087 9367
rect 3617 9333 3651 9367
rect 4353 9333 4387 9367
rect 4537 9333 4571 9367
rect 7757 9333 7791 9367
rect 9781 9333 9815 9367
rect 11529 9333 11563 9367
rect 13185 9333 13219 9367
rect 15301 9333 15335 9367
rect 15485 9333 15519 9367
rect 15761 9333 15795 9367
rect 17325 9333 17359 9367
rect 17509 9333 17543 9367
rect 17785 9333 17819 9367
rect 17969 9333 18003 9367
rect 18429 9333 18463 9367
rect 21005 9333 21039 9367
rect 21189 9333 21223 9367
rect 21833 9333 21867 9367
rect 2053 9129 2087 9163
rect 2513 9129 2547 9163
rect 2881 9129 2915 9163
rect 3525 9129 3559 9163
rect 4261 9129 4295 9163
rect 6561 9129 6595 9163
rect 6837 9129 6871 9163
rect 7021 9129 7055 9163
rect 11253 9129 11287 9163
rect 11805 9129 11839 9163
rect 12081 9129 12115 9163
rect 13553 9129 13587 9163
rect 14105 9129 14139 9163
rect 14473 9129 14507 9163
rect 16635 9129 16669 9163
rect 18337 9129 18371 9163
rect 18613 9129 18647 9163
rect 22293 9129 22327 9163
rect 22569 9129 22603 9163
rect 4169 9061 4203 9095
rect 4813 9061 4847 9095
rect 5365 9061 5399 9095
rect 18153 9061 18187 9095
rect 5089 8993 5123 9027
rect 6009 8993 6043 9027
rect 6193 8993 6227 9027
rect 9873 8993 9907 9027
rect 14841 8993 14875 9027
rect 20545 8993 20579 9027
rect 2237 8925 2271 8959
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 3433 8925 3467 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 5273 8925 5307 8959
rect 5716 8925 5750 8959
rect 5825 8925 5859 8959
rect 6101 8925 6135 8959
rect 6377 8925 6411 8959
rect 9597 8925 9631 8959
rect 9689 8925 9723 8959
rect 11529 8925 11563 8959
rect 12265 8925 12299 8959
rect 12357 8925 12391 8959
rect 12541 8925 12575 8959
rect 12633 8925 12667 8959
rect 13001 8925 13035 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 14565 8925 14599 8959
rect 15209 8925 15243 8959
rect 18061 8925 18095 8959
rect 18245 8925 18279 8959
rect 18521 8925 18555 8959
rect 18613 8925 18647 8959
rect 18797 8925 18831 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 20269 8925 20303 8959
rect 22477 8925 22511 8959
rect 24409 8925 24443 8959
rect 2329 8857 2363 8891
rect 2529 8857 2563 8891
rect 3249 8857 3283 8891
rect 3801 8857 3835 8891
rect 6653 8857 6687 8891
rect 6853 8857 6887 8891
rect 10140 8857 10174 8891
rect 13185 8857 13219 8891
rect 13277 8857 13311 8891
rect 17785 8857 17819 8891
rect 20361 8857 20395 8891
rect 20821 8857 20855 8891
rect 2697 8789 2731 8823
rect 5549 8789 5583 8823
rect 11989 8789 12023 8823
rect 18981 8789 19015 8823
rect 19349 8789 19383 8823
rect 24501 8789 24535 8823
rect 1593 8585 1627 8619
rect 5273 8585 5307 8619
rect 9505 8585 9539 8619
rect 12541 8585 12575 8619
rect 16313 8585 16347 8619
rect 17877 8585 17911 8619
rect 22477 8585 22511 8619
rect 22661 8585 22695 8619
rect 25145 8585 25179 8619
rect 3801 8517 3835 8551
rect 4017 8517 4051 8551
rect 4721 8517 4755 8551
rect 12909 8517 12943 8551
rect 16129 8517 16163 8551
rect 16681 8517 16715 8551
rect 23673 8517 23707 8551
rect 1409 8449 1443 8483
rect 5457 8449 5491 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 5917 8449 5951 8483
rect 8125 8449 8159 8483
rect 8392 8449 8426 8483
rect 11529 8449 11563 8483
rect 12081 8449 12115 8483
rect 13093 8449 13127 8483
rect 13185 8449 13219 8483
rect 13461 8449 13495 8483
rect 13553 8449 13587 8483
rect 13921 8449 13955 8483
rect 15761 8449 15795 8483
rect 16957 8449 16991 8483
rect 18153 8449 18187 8483
rect 18429 8449 18463 8483
rect 18613 8449 18647 8483
rect 22569 8449 22603 8483
rect 23397 8449 23431 8483
rect 25605 8449 25639 8483
rect 5181 8381 5215 8415
rect 16773 8381 16807 8415
rect 21925 8381 21959 8415
rect 5089 8313 5123 8347
rect 11989 8313 12023 8347
rect 14105 8313 14139 8347
rect 18245 8313 18279 8347
rect 25881 8313 25915 8347
rect 3985 8245 4019 8279
rect 4169 8245 4203 8279
rect 11805 8245 11839 8279
rect 12173 8245 12207 8279
rect 13369 8245 13403 8279
rect 13921 8245 13955 8279
rect 16129 8245 16163 8279
rect 16681 8245 16715 8279
rect 17141 8245 17175 8279
rect 18337 8245 18371 8279
rect 3433 8041 3467 8075
rect 4537 8041 4571 8075
rect 5917 8041 5951 8075
rect 6285 8041 6319 8075
rect 7941 8041 7975 8075
rect 9689 8041 9723 8075
rect 13001 8041 13035 8075
rect 13737 8041 13771 8075
rect 13921 8041 13955 8075
rect 15393 8041 15427 8075
rect 15577 8041 15611 8075
rect 16957 8041 16991 8075
rect 17877 8041 17911 8075
rect 18061 8041 18095 8075
rect 18521 8041 18555 8075
rect 19717 8041 19751 8075
rect 3065 7973 3099 8007
rect 3801 7973 3835 8007
rect 4721 7973 4755 8007
rect 5641 7973 5675 8007
rect 15025 7973 15059 8007
rect 18705 7973 18739 8007
rect 19533 7973 19567 8007
rect 2697 7905 2731 7939
rect 5733 7905 5767 7939
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 5273 7837 5307 7871
rect 5825 7837 5859 7871
rect 8125 7837 8159 7871
rect 9965 7837 9999 7871
rect 10241 7837 10275 7871
rect 10425 7837 10459 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 13461 7837 13495 7871
rect 17509 7837 17543 7871
rect 18153 7837 18187 7871
rect 22661 7837 22695 7871
rect 3249 7769 3283 7803
rect 4353 7769 4387 7803
rect 4569 7769 4603 7803
rect 9689 7769 9723 7803
rect 13553 7769 13587 7803
rect 15669 7769 15703 7803
rect 19257 7769 19291 7803
rect 3157 7701 3191 7735
rect 3449 7701 3483 7735
rect 3617 7701 3651 7735
rect 9873 7701 9907 7735
rect 10333 7701 10367 7735
rect 13753 7701 13787 7735
rect 15393 7701 15427 7735
rect 17877 7701 17911 7735
rect 18521 7701 18555 7735
rect 23213 7701 23247 7735
rect 2329 7497 2363 7531
rect 3985 7497 4019 7531
rect 10057 7497 10091 7531
rect 11713 7497 11747 7531
rect 12081 7497 12115 7531
rect 18613 7497 18647 7531
rect 19165 7497 19199 7531
rect 23627 7497 23661 7531
rect 2850 7429 2884 7463
rect 10885 7429 10919 7463
rect 11085 7429 11119 7463
rect 18429 7429 18463 7463
rect 18705 7429 18739 7463
rect 24041 7429 24075 7463
rect 2513 7361 2547 7395
rect 4261 7361 4295 7395
rect 4905 7361 4939 7395
rect 8217 7361 8251 7395
rect 8484 7361 8518 7395
rect 9781 7361 9815 7395
rect 9873 7361 9907 7395
rect 10793 7361 10827 7395
rect 11529 7361 11563 7395
rect 11897 7361 11931 7395
rect 18061 7361 18095 7395
rect 20729 7361 20763 7395
rect 21465 7361 21499 7395
rect 21833 7361 21867 7395
rect 23765 7361 23799 7395
rect 2605 7293 2639 7327
rect 4353 7293 4387 7327
rect 10241 7293 10275 7327
rect 20545 7293 20579 7327
rect 20637 7293 20671 7327
rect 20821 7293 20855 7327
rect 21557 7293 21591 7327
rect 22201 7293 22235 7327
rect 4629 7225 4663 7259
rect 19073 7225 19107 7259
rect 4721 7157 4755 7191
rect 9597 7157 9631 7191
rect 11069 7157 11103 7191
rect 11253 7157 11287 7191
rect 18429 7157 18463 7191
rect 20361 7157 20395 7191
rect 5181 6953 5215 6987
rect 6101 6953 6135 6987
rect 6469 6953 6503 6987
rect 7481 6953 7515 6987
rect 7665 6953 7699 6987
rect 9137 6953 9171 6987
rect 9505 6953 9539 6987
rect 10793 6953 10827 6987
rect 15163 6953 15197 6987
rect 18291 6953 18325 6987
rect 18889 6953 18923 6987
rect 21143 6953 21177 6987
rect 8677 6885 8711 6919
rect 15301 6885 15335 6919
rect 18751 6885 18785 6919
rect 6285 6817 6319 6851
rect 9597 6817 9631 6851
rect 10885 6817 10919 6851
rect 16497 6817 16531 6851
rect 19349 6817 19383 6851
rect 22385 6817 22419 6851
rect 3801 6749 3835 6783
rect 5825 6749 5859 6783
rect 6377 6749 6411 6783
rect 6929 6749 6963 6783
rect 8309 6749 8343 6783
rect 9045 6749 9079 6783
rect 11069 6749 11103 6783
rect 12633 6749 12667 6783
rect 13645 6749 13679 6783
rect 14381 6749 14415 6783
rect 15025 6749 15059 6783
rect 15485 6749 15519 6783
rect 15669 6749 15703 6783
rect 16037 6749 16071 6783
rect 16865 6749 16899 6783
rect 18613 6749 18647 6783
rect 19073 6749 19107 6783
rect 19717 6749 19751 6783
rect 21281 6749 21315 6783
rect 22293 6749 22327 6783
rect 23765 6749 23799 6783
rect 24041 6749 24075 6783
rect 4068 6681 4102 6715
rect 7297 6681 7331 6715
rect 10517 6681 10551 6715
rect 10977 6681 11011 6715
rect 11336 6681 11370 6715
rect 14933 6681 14967 6715
rect 15853 6681 15887 6715
rect 15945 6681 15979 6715
rect 21373 6681 21407 6715
rect 6837 6613 6871 6647
rect 7021 6613 7055 6647
rect 7507 6613 7541 6647
rect 8769 6613 8803 6647
rect 10241 6613 10275 6647
rect 10609 6613 10643 6647
rect 12449 6613 12483 6647
rect 13185 6613 13219 6647
rect 13737 6613 13771 6647
rect 15393 6613 15427 6647
rect 16221 6613 16255 6647
rect 19073 6613 19107 6647
rect 23857 6613 23891 6647
rect 24133 6613 24167 6647
rect 6377 6409 6411 6443
rect 8953 6409 8987 6443
rect 9137 6409 9171 6443
rect 10333 6409 10367 6443
rect 12173 6409 12207 6443
rect 15117 6409 15151 6443
rect 17601 6409 17635 6443
rect 20729 6409 20763 6443
rect 22759 6409 22793 6443
rect 4997 6341 5031 6375
rect 5825 6341 5859 6375
rect 5917 6341 5951 6375
rect 6745 6341 6779 6375
rect 8401 6341 8435 6375
rect 11345 6341 11379 6375
rect 12265 6341 12299 6375
rect 12725 6341 12759 6375
rect 15209 6341 15243 6375
rect 20361 6341 20395 6375
rect 20821 6341 20855 6375
rect 5549 6273 5583 6307
rect 5697 6273 5731 6307
rect 6055 6273 6089 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 6929 6273 6963 6307
rect 7021 6273 7055 6307
rect 7849 6273 7883 6307
rect 9134 6273 9168 6307
rect 9689 6273 9723 6307
rect 9837 6273 9871 6307
rect 9965 6273 9999 6307
rect 10057 6273 10091 6307
rect 10195 6273 10229 6307
rect 10425 6273 10459 6307
rect 11529 6273 11563 6307
rect 12449 6273 12483 6307
rect 12909 6273 12943 6307
rect 13277 6273 13311 6307
rect 14933 6273 14967 6307
rect 15117 6273 15151 6307
rect 15485 6273 15519 6307
rect 16037 6273 16071 6307
rect 16221 6273 16255 6307
rect 16314 6273 16348 6307
rect 16865 6273 16899 6307
rect 17141 6273 17175 6307
rect 17509 6273 17543 6307
rect 19257 6273 19291 6307
rect 19441 6273 19475 6307
rect 19533 6273 19567 6307
rect 19717 6273 19751 6307
rect 19809 6273 19843 6307
rect 20177 6273 20211 6307
rect 20453 6273 20487 6307
rect 20545 6273 20579 6307
rect 21005 6273 21039 6307
rect 21189 6273 21223 6307
rect 21281 6273 21315 6307
rect 21833 6273 21867 6307
rect 22017 6273 22051 6307
rect 22293 6273 22327 6307
rect 22477 6273 22511 6307
rect 22661 6273 22695 6307
rect 22845 6273 22879 6307
rect 22937 6273 22971 6307
rect 23397 6273 23431 6307
rect 5457 6205 5491 6239
rect 7113 6205 7147 6239
rect 7573 6205 7607 6239
rect 9597 6205 9631 6239
rect 10517 6205 10551 6239
rect 10793 6205 10827 6239
rect 12633 6205 12667 6239
rect 15301 6205 15335 6239
rect 16129 6205 16163 6239
rect 17049 6205 17083 6239
rect 23029 6205 23063 6239
rect 5365 6137 5399 6171
rect 6193 6137 6227 6171
rect 7389 6137 7423 6171
rect 8677 6137 8711 6171
rect 9505 6137 9539 6171
rect 16957 6137 16991 6171
rect 19349 6137 19383 6171
rect 7941 6069 7975 6103
rect 8309 6069 8343 6103
rect 8861 6069 8895 6103
rect 12541 6069 12575 6103
rect 14703 6069 14737 6103
rect 15209 6069 15243 6103
rect 15669 6069 15703 6103
rect 15853 6069 15887 6103
rect 16681 6069 16715 6103
rect 19717 6069 19751 6103
rect 19993 6069 20027 6103
rect 22201 6069 22235 6103
rect 22293 6069 22327 6103
rect 24823 6069 24857 6103
rect 6745 5865 6779 5899
rect 9781 5865 9815 5899
rect 10057 5865 10091 5899
rect 12817 5865 12851 5899
rect 14197 5865 14231 5899
rect 14749 5865 14783 5899
rect 15025 5865 15059 5899
rect 17693 5865 17727 5899
rect 20453 5865 20487 5899
rect 20913 5865 20947 5899
rect 22293 5865 22327 5899
rect 7481 5797 7515 5831
rect 7573 5797 7607 5831
rect 8585 5797 8619 5831
rect 10793 5797 10827 5831
rect 11345 5797 11379 5831
rect 17877 5797 17911 5831
rect 25053 5797 25087 5831
rect 7113 5729 7147 5763
rect 7665 5729 7699 5763
rect 8309 5729 8343 5763
rect 8769 5729 8803 5763
rect 10517 5729 10551 5763
rect 17417 5729 17451 5763
rect 22385 5729 22419 5763
rect 5273 5661 5307 5695
rect 7849 5661 7883 5695
rect 9137 5661 9171 5695
rect 9230 5661 9264 5695
rect 9602 5661 9636 5695
rect 10241 5661 10275 5695
rect 10333 5661 10367 5695
rect 10609 5661 10643 5695
rect 11437 5661 11471 5695
rect 14105 5661 14139 5695
rect 15209 5661 15243 5695
rect 15485 5661 15519 5695
rect 15669 5661 15703 5695
rect 17969 5661 18003 5695
rect 20361 5661 20395 5695
rect 22109 5661 22143 5695
rect 22753 5661 22787 5695
rect 24869 5661 24903 5695
rect 9413 5593 9447 5627
rect 9505 5593 9539 5627
rect 10977 5593 11011 5627
rect 11704 5593 11738 5627
rect 14565 5593 14599 5627
rect 17509 5593 17543 5627
rect 20729 5593 20763 5627
rect 20945 5593 20979 5627
rect 21925 5593 21959 5627
rect 8033 5525 8067 5559
rect 11069 5525 11103 5559
rect 11161 5525 11195 5559
rect 14765 5525 14799 5559
rect 14933 5525 14967 5559
rect 15393 5525 15427 5559
rect 17709 5525 17743 5559
rect 18061 5525 18095 5559
rect 21097 5525 21131 5559
rect 24179 5525 24213 5559
rect 6377 5321 6411 5355
rect 7221 5321 7255 5355
rect 7665 5321 7699 5355
rect 10241 5321 10275 5355
rect 15577 5321 15611 5355
rect 16405 5321 16439 5355
rect 16773 5321 16807 5355
rect 20290 5321 20324 5355
rect 20453 5321 20487 5355
rect 22385 5321 22419 5355
rect 7021 5253 7055 5287
rect 19349 5253 19383 5287
rect 19549 5253 19583 5287
rect 20085 5253 20119 5287
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 6929 5185 6963 5219
rect 7481 5185 7515 5219
rect 7665 5185 7699 5219
rect 7757 5185 7791 5219
rect 7849 5185 7883 5219
rect 10425 5185 10459 5219
rect 14289 5185 14323 5219
rect 15761 5185 15795 5219
rect 16313 5185 16347 5219
rect 16957 5185 16991 5219
rect 17049 5185 17083 5219
rect 17233 5185 17267 5219
rect 17417 5185 17451 5219
rect 22293 5185 22327 5219
rect 22477 5185 22511 5219
rect 22661 5185 22695 5219
rect 22845 5185 22879 5219
rect 22937 5185 22971 5219
rect 6837 5117 6871 5151
rect 10701 5117 10735 5151
rect 14105 5117 14139 5151
rect 15853 5117 15887 5151
rect 15945 5117 15979 5151
rect 16037 5117 16071 5151
rect 17693 5117 17727 5151
rect 7389 5049 7423 5083
rect 17141 5049 17175 5083
rect 22661 5049 22695 5083
rect 7205 4981 7239 5015
rect 10609 4981 10643 5015
rect 14473 4981 14507 5015
rect 17509 4981 17543 5015
rect 17969 4981 18003 5015
rect 19533 4981 19567 5015
rect 19717 4981 19751 5015
rect 20269 4981 20303 5015
rect 6193 4777 6227 4811
rect 10977 4777 11011 4811
rect 12081 4777 12115 4811
rect 25973 4777 26007 4811
rect 6377 4709 6411 4743
rect 13553 4709 13587 4743
rect 18981 4709 19015 4743
rect 20177 4709 20211 4743
rect 14933 4641 14967 4675
rect 19533 4641 19567 4675
rect 19625 4641 19659 4675
rect 20269 4641 20303 4675
rect 20545 4641 20579 4675
rect 20821 4641 20855 4675
rect 21281 4641 21315 4675
rect 21741 4641 21775 4675
rect 22017 4641 22051 4675
rect 5181 4573 5215 4607
rect 5641 4573 5675 4607
rect 5917 4573 5951 4607
rect 6469 4573 6503 4607
rect 7665 4573 7699 4607
rect 7849 4573 7883 4607
rect 8493 4573 8527 4607
rect 10885 4573 10919 4607
rect 11069 4573 11103 4607
rect 11161 4573 11195 4607
rect 11345 4573 11379 4607
rect 11989 4573 12023 4607
rect 13737 4573 13771 4607
rect 13829 4573 13863 4607
rect 14289 4573 14323 4607
rect 14467 4573 14501 4607
rect 15209 4573 15243 4607
rect 16589 4573 16623 4607
rect 16773 4573 16807 4607
rect 18889 4573 18923 4607
rect 19441 4573 19475 4607
rect 19717 4573 19751 4607
rect 19901 4573 19935 4607
rect 20085 4573 20119 4607
rect 20361 4573 20395 4607
rect 20729 4573 20763 4607
rect 20913 4573 20947 4607
rect 21005 4573 21039 4607
rect 21189 4573 21223 4607
rect 21649 4573 21683 4607
rect 22109 4573 22143 4607
rect 22293 4573 22327 4607
rect 25789 4573 25823 4607
rect 5457 4505 5491 4539
rect 6009 4505 6043 4539
rect 11253 4505 11287 4539
rect 13553 4505 13587 4539
rect 14381 4505 14415 4539
rect 14565 4505 14599 4539
rect 14749 4505 14783 4539
rect 15025 4505 15059 4539
rect 4997 4437 5031 4471
rect 5825 4437 5859 4471
rect 6209 4437 6243 4471
rect 6561 4437 6595 4471
rect 7757 4437 7791 4471
rect 8309 4437 8343 4471
rect 15393 4437 15427 4471
rect 16957 4437 16991 4471
rect 19257 4437 19291 4471
rect 22477 4437 22511 4471
rect 5733 4233 5767 4267
rect 7865 4233 7899 4267
rect 9505 4233 9539 4267
rect 11253 4233 11287 4267
rect 11897 4233 11931 4267
rect 13369 4233 13403 4267
rect 20085 4233 20119 4267
rect 4620 4165 4654 4199
rect 5825 4165 5859 4199
rect 6041 4165 6075 4199
rect 7021 4165 7055 4199
rect 7221 4165 7255 4199
rect 7665 4165 7699 4199
rect 10057 4165 10091 4199
rect 11529 4165 11563 4199
rect 11713 4165 11747 4199
rect 16957 4165 16991 4199
rect 22845 4165 22879 4199
rect 22937 4165 22971 4199
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 6929 4097 6963 4131
rect 8125 4097 8159 4131
rect 8392 4097 8426 4131
rect 10241 4097 10275 4131
rect 10333 4097 10367 4131
rect 10609 4097 10643 4131
rect 11069 4097 11103 4131
rect 11345 4097 11379 4131
rect 11989 4097 12023 4131
rect 12633 4097 12667 4131
rect 12909 4097 12943 4131
rect 13185 4097 13219 4131
rect 14105 4097 14139 4131
rect 14565 4097 14599 4131
rect 14749 4097 14783 4131
rect 15025 4097 15059 4131
rect 16129 4097 16163 4131
rect 16865 4097 16899 4131
rect 17049 4097 17083 4131
rect 17167 4097 17201 4131
rect 18337 4097 18371 4131
rect 20453 4097 20487 4131
rect 20821 4097 20855 4131
rect 21097 4097 21131 4131
rect 22201 4097 22235 4131
rect 22661 4097 22695 4131
rect 23029 4097 23063 4131
rect 4353 4029 4387 4063
rect 10701 4029 10735 4063
rect 14197 4029 14231 4063
rect 14473 4029 14507 4063
rect 16221 4029 16255 4063
rect 17325 4029 17359 4063
rect 18613 4029 18647 4063
rect 20361 4029 20395 4063
rect 20729 4029 20763 4063
rect 21005 4029 21039 4063
rect 22293 4029 22327 4063
rect 22569 4029 22603 4063
rect 7389 3961 7423 3995
rect 10977 3961 11011 3995
rect 15577 3961 15611 3995
rect 16497 3961 16531 3995
rect 20177 3961 20211 3995
rect 21465 3961 21499 3995
rect 6009 3893 6043 3927
rect 6193 3893 6227 3927
rect 6469 3893 6503 3927
rect 7205 3893 7239 3927
rect 7849 3893 7883 3927
rect 8033 3893 8067 3927
rect 10057 3893 10091 3927
rect 11069 3893 11103 3927
rect 13001 3893 13035 3927
rect 14565 3893 14599 3927
rect 16681 3893 16715 3927
rect 23213 3893 23247 3927
rect 7297 3689 7331 3723
rect 8493 3689 8527 3723
rect 11805 3689 11839 3723
rect 14749 3689 14783 3723
rect 17601 3689 17635 3723
rect 21005 3689 21039 3723
rect 22937 3689 22971 3723
rect 23581 3689 23615 3723
rect 7021 3621 7055 3655
rect 8677 3621 8711 3655
rect 13875 3621 13909 3655
rect 15761 3621 15795 3655
rect 5273 3553 5307 3587
rect 7941 3553 7975 3587
rect 8217 3553 8251 3587
rect 8953 3553 8987 3587
rect 12081 3553 12115 3587
rect 14381 3553 14415 3587
rect 14657 3553 14691 3587
rect 15853 3553 15887 3587
rect 19257 3553 19291 3587
rect 21189 3553 21223 3587
rect 21557 3553 21591 3587
rect 4905 3485 4939 3519
rect 5181 3485 5215 3519
rect 5641 3485 5675 3519
rect 7849 3485 7883 3519
rect 10425 3485 10459 3519
rect 10692 3485 10726 3519
rect 12449 3485 12483 3519
rect 14289 3485 14323 3519
rect 14749 3485 14783 3519
rect 15025 3485 15059 3519
rect 15209 3485 15243 3519
rect 15393 3485 15427 3519
rect 15577 3485 15611 3519
rect 16221 3485 16255 3519
rect 17785 3485 17819 3519
rect 18061 3485 18095 3519
rect 18889 3485 18923 3519
rect 18981 3485 19015 3519
rect 19625 3485 19659 3519
rect 23397 3485 23431 3519
rect 5908 3417 5942 3451
rect 7113 3417 7147 3451
rect 8309 3417 8343 3451
rect 8509 3417 8543 3451
rect 9198 3417 9232 3451
rect 15485 3417 15519 3451
rect 4721 3349 4755 3383
rect 5549 3349 5583 3383
rect 7313 3349 7347 3383
rect 7481 3349 7515 3383
rect 10333 3349 10367 3383
rect 14933 3349 14967 3383
rect 17877 3349 17911 3383
rect 18153 3349 18187 3383
rect 6101 3145 6135 3179
rect 6837 3145 6871 3179
rect 8493 3145 8527 3179
rect 11345 3145 11379 3179
rect 14519 3145 14553 3179
rect 16405 3145 16439 3179
rect 20269 3145 20303 3179
rect 20453 3145 20487 3179
rect 21373 3145 21407 3179
rect 6377 3077 6411 3111
rect 10210 3077 10244 3111
rect 18521 3077 18555 3111
rect 4721 3009 4755 3043
rect 4977 3009 5011 3043
rect 8677 3009 8711 3043
rect 9965 3009 9999 3043
rect 13093 3009 13127 3043
rect 16313 3009 16347 3043
rect 16681 3009 16715 3043
rect 19441 3009 19475 3043
rect 19993 3009 20027 3043
rect 20361 3009 20395 3043
rect 21281 3009 21315 3043
rect 12725 2941 12759 2975
rect 17049 2941 17083 2975
rect 19717 2941 19751 2975
rect 20269 2941 20303 2975
rect 6653 2873 6687 2907
rect 20085 2873 20119 2907
rect 6009 2601 6043 2635
rect 8033 2601 8067 2635
rect 11897 2601 11931 2635
rect 13829 2601 13863 2635
rect 15577 2601 15611 2635
rect 23949 2601 23983 2635
rect 1501 2397 1535 2431
rect 3985 2397 4019 2431
rect 6193 2397 6227 2431
rect 7849 2397 7883 2431
rect 11713 2397 11747 2431
rect 13737 2397 13771 2431
rect 15761 2397 15795 2431
rect 20177 2397 20211 2431
rect 24133 2397 24167 2431
rect 1869 2329 1903 2363
rect 25605 2329 25639 2363
rect 4169 2261 4203 2295
rect 20269 2261 20303 2295
rect 25697 2261 25731 2295
<< metal1 >>
rect 1104 27226 26312 27248
rect 1104 27174 4761 27226
rect 4813 27174 4825 27226
rect 4877 27174 4889 27226
rect 4941 27174 4953 27226
rect 5005 27174 5017 27226
rect 5069 27174 11063 27226
rect 11115 27174 11127 27226
rect 11179 27174 11191 27226
rect 11243 27174 11255 27226
rect 11307 27174 11319 27226
rect 11371 27174 17365 27226
rect 17417 27174 17429 27226
rect 17481 27174 17493 27226
rect 17545 27174 17557 27226
rect 17609 27174 17621 27226
rect 17673 27174 23667 27226
rect 23719 27174 23731 27226
rect 23783 27174 23795 27226
rect 23847 27174 23859 27226
rect 23911 27174 23923 27226
rect 23975 27174 26312 27226
rect 1104 27152 26312 27174
rect 3234 27072 3240 27124
rect 3292 27112 3298 27124
rect 3973 27115 4031 27121
rect 3973 27112 3985 27115
rect 3292 27084 3985 27112
rect 3292 27072 3298 27084
rect 3973 27081 3985 27084
rect 4019 27081 4031 27115
rect 3973 27075 4031 27081
rect 7098 27072 7104 27124
rect 7156 27112 7162 27124
rect 7377 27115 7435 27121
rect 7377 27112 7389 27115
rect 7156 27084 7389 27112
rect 7156 27072 7162 27084
rect 7377 27081 7389 27084
rect 7423 27081 7435 27115
rect 7377 27075 7435 27081
rect 11606 27072 11612 27124
rect 11664 27112 11670 27124
rect 12069 27115 12127 27121
rect 12069 27112 12081 27115
rect 11664 27084 12081 27112
rect 11664 27072 11670 27084
rect 12069 27081 12081 27084
rect 12115 27081 12127 27115
rect 12069 27075 12127 27081
rect 19334 27072 19340 27124
rect 19392 27112 19398 27124
rect 19613 27115 19671 27121
rect 19613 27112 19625 27115
rect 19392 27084 19625 27112
rect 19392 27072 19398 27084
rect 19613 27081 19625 27084
rect 19659 27081 19671 27115
rect 19613 27075 19671 27081
rect 23474 27072 23480 27124
rect 23532 27072 23538 27124
rect 3881 27047 3939 27053
rect 3881 27013 3893 27047
rect 3927 27044 3939 27047
rect 10778 27044 10784 27056
rect 3927 27016 10784 27044
rect 3927 27013 3939 27016
rect 3881 27007 3939 27013
rect 10778 27004 10784 27016
rect 10836 27004 10842 27056
rect 1394 26936 1400 26988
rect 1452 26936 1458 26988
rect 7285 26979 7343 26985
rect 7285 26945 7297 26979
rect 7331 26976 7343 26979
rect 11514 26976 11520 26988
rect 7331 26948 11520 26976
rect 7331 26945 7343 26948
rect 7285 26939 7343 26945
rect 11514 26936 11520 26948
rect 11572 26936 11578 26988
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12342 26976 12348 26988
rect 11931 26948 12348 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12342 26936 12348 26948
rect 12400 26936 12406 26988
rect 15470 26936 15476 26988
rect 15528 26976 15534 26988
rect 15749 26979 15807 26985
rect 15749 26976 15761 26979
rect 15528 26948 15761 26976
rect 15528 26936 15534 26948
rect 15749 26945 15761 26948
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 19334 26936 19340 26988
rect 19392 26976 19398 26988
rect 19521 26979 19579 26985
rect 19521 26976 19533 26979
rect 19392 26948 19533 26976
rect 19392 26936 19398 26948
rect 19521 26945 19533 26948
rect 19567 26945 19579 26979
rect 19521 26939 19579 26945
rect 23382 26936 23388 26988
rect 23440 26936 23446 26988
rect 1581 26775 1639 26781
rect 1581 26741 1593 26775
rect 1627 26772 1639 26775
rect 2590 26772 2596 26784
rect 1627 26744 2596 26772
rect 1627 26741 1639 26744
rect 1581 26735 1639 26741
rect 2590 26732 2596 26744
rect 2648 26732 2654 26784
rect 15565 26775 15623 26781
rect 15565 26741 15577 26775
rect 15611 26772 15623 26775
rect 16298 26772 16304 26784
rect 15611 26744 16304 26772
rect 15611 26741 15623 26744
rect 15565 26735 15623 26741
rect 16298 26732 16304 26744
rect 16356 26732 16362 26784
rect 1104 26682 26312 26704
rect 1104 26630 4101 26682
rect 4153 26630 4165 26682
rect 4217 26630 4229 26682
rect 4281 26630 4293 26682
rect 4345 26630 4357 26682
rect 4409 26630 10403 26682
rect 10455 26630 10467 26682
rect 10519 26630 10531 26682
rect 10583 26630 10595 26682
rect 10647 26630 10659 26682
rect 10711 26630 16705 26682
rect 16757 26630 16769 26682
rect 16821 26630 16833 26682
rect 16885 26630 16897 26682
rect 16949 26630 16961 26682
rect 17013 26630 23007 26682
rect 23059 26630 23071 26682
rect 23123 26630 23135 26682
rect 23187 26630 23199 26682
rect 23251 26630 23263 26682
rect 23315 26630 26312 26682
rect 1104 26608 26312 26630
rect 9674 26460 9680 26512
rect 9732 26460 9738 26512
rect 15672 26472 19104 26500
rect 6825 26435 6883 26441
rect 6825 26401 6837 26435
rect 6871 26432 6883 26435
rect 9858 26432 9864 26444
rect 6871 26404 9864 26432
rect 6871 26401 6883 26404
rect 6825 26395 6883 26401
rect 9858 26392 9864 26404
rect 9916 26392 9922 26444
rect 13722 26392 13728 26444
rect 13780 26432 13786 26444
rect 13780 26404 15332 26432
rect 13780 26392 13786 26404
rect 6546 26324 6552 26376
rect 6604 26324 6610 26376
rect 8938 26324 8944 26376
rect 8996 26364 9002 26376
rect 8996 26336 9904 26364
rect 8996 26324 9002 26336
rect 7466 26256 7472 26308
rect 7524 26256 7530 26308
rect 9214 26256 9220 26308
rect 9272 26256 9278 26308
rect 9398 26256 9404 26308
rect 9456 26256 9462 26308
rect 9876 26305 9904 26336
rect 9950 26324 9956 26376
rect 10008 26324 10014 26376
rect 11882 26324 11888 26376
rect 11940 26364 11946 26376
rect 12069 26367 12127 26373
rect 12069 26364 12081 26367
rect 11940 26336 12081 26364
rect 11940 26324 11946 26336
rect 12069 26333 12081 26336
rect 12115 26333 12127 26367
rect 12069 26327 12127 26333
rect 12434 26324 12440 26376
rect 12492 26324 12498 26376
rect 13814 26324 13820 26376
rect 13872 26324 13878 26376
rect 15304 26373 15332 26404
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26364 15347 26367
rect 15672 26364 15700 26472
rect 16301 26435 16359 26441
rect 16301 26401 16313 26435
rect 16347 26432 16359 26435
rect 17313 26435 17371 26441
rect 17313 26432 17325 26435
rect 16347 26404 17325 26432
rect 16347 26401 16359 26404
rect 16301 26395 16359 26401
rect 17313 26401 17325 26404
rect 17359 26401 17371 26435
rect 17313 26395 17371 26401
rect 17497 26435 17555 26441
rect 17497 26401 17509 26435
rect 17543 26432 17555 26435
rect 18414 26432 18420 26444
rect 17543 26404 18420 26432
rect 17543 26401 17555 26404
rect 17497 26395 17555 26401
rect 18414 26392 18420 26404
rect 18472 26392 18478 26444
rect 19076 26376 19104 26472
rect 20257 26435 20315 26441
rect 20257 26401 20269 26435
rect 20303 26432 20315 26435
rect 20714 26432 20720 26444
rect 20303 26404 20720 26432
rect 20303 26401 20315 26404
rect 20257 26395 20315 26401
rect 20714 26392 20720 26404
rect 20772 26392 20778 26444
rect 15335 26336 15700 26364
rect 15749 26367 15807 26373
rect 15335 26333 15347 26336
rect 15289 26327 15347 26333
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 15930 26364 15936 26376
rect 15795 26336 15936 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 15930 26324 15936 26336
rect 15988 26324 15994 26376
rect 16574 26324 16580 26376
rect 16632 26364 16638 26376
rect 17221 26367 17279 26373
rect 17221 26364 17233 26367
rect 16632 26336 17233 26364
rect 16632 26324 16638 26336
rect 17221 26333 17233 26336
rect 17267 26333 17279 26367
rect 17221 26327 17279 26333
rect 9677 26299 9735 26305
rect 9677 26265 9689 26299
rect 9723 26265 9735 26299
rect 9677 26259 9735 26265
rect 9861 26299 9919 26305
rect 9861 26265 9873 26299
rect 9907 26296 9919 26299
rect 10594 26296 10600 26308
rect 9907 26268 10600 26296
rect 9907 26265 9919 26268
rect 9861 26259 9919 26265
rect 8294 26188 8300 26240
rect 8352 26188 8358 26240
rect 9582 26188 9588 26240
rect 9640 26188 9646 26240
rect 9692 26228 9720 26259
rect 10594 26256 10600 26268
rect 10652 26256 10658 26308
rect 13832 26296 13860 26324
rect 13478 26268 13860 26296
rect 15381 26299 15439 26305
rect 15381 26265 15393 26299
rect 15427 26296 15439 26299
rect 15470 26296 15476 26308
rect 15427 26268 15476 26296
rect 15427 26265 15439 26268
rect 15381 26259 15439 26265
rect 15470 26256 15476 26268
rect 15528 26256 15534 26308
rect 17236 26296 17264 26327
rect 17402 26324 17408 26376
rect 17460 26324 17466 26376
rect 17770 26324 17776 26376
rect 17828 26364 17834 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 17828 26336 18061 26364
rect 17828 26324 17834 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 18049 26327 18107 26333
rect 19058 26324 19064 26376
rect 19116 26364 19122 26376
rect 20165 26367 20223 26373
rect 20165 26364 20177 26367
rect 19116 26336 20177 26364
rect 19116 26324 19122 26336
rect 20165 26333 20177 26336
rect 20211 26364 20223 26367
rect 20441 26367 20499 26373
rect 20441 26364 20453 26367
rect 20211 26336 20453 26364
rect 20211 26333 20223 26336
rect 20165 26327 20223 26333
rect 20441 26333 20453 26336
rect 20487 26333 20499 26367
rect 20441 26327 20499 26333
rect 17681 26299 17739 26305
rect 17681 26296 17693 26299
rect 17236 26268 17693 26296
rect 17681 26265 17693 26268
rect 17727 26265 17739 26299
rect 17681 26259 17739 26265
rect 17865 26299 17923 26305
rect 17865 26265 17877 26299
rect 17911 26265 17923 26299
rect 17865 26259 17923 26265
rect 20533 26299 20591 26305
rect 20533 26265 20545 26299
rect 20579 26296 20591 26299
rect 20806 26296 20812 26308
rect 20579 26268 20812 26296
rect 20579 26265 20591 26268
rect 20533 26259 20591 26265
rect 9766 26228 9772 26240
rect 9692 26200 9772 26228
rect 9766 26188 9772 26200
rect 9824 26228 9830 26240
rect 10870 26228 10876 26240
rect 9824 26200 10876 26228
rect 9824 26188 9830 26200
rect 10870 26188 10876 26200
rect 10928 26188 10934 26240
rect 13863 26231 13921 26237
rect 13863 26197 13875 26231
rect 13909 26228 13921 26231
rect 14642 26228 14648 26240
rect 13909 26200 14648 26228
rect 13909 26197 13921 26200
rect 13863 26191 13921 26197
rect 14642 26188 14648 26200
rect 14700 26188 14706 26240
rect 17037 26231 17095 26237
rect 17037 26197 17049 26231
rect 17083 26228 17095 26231
rect 17218 26228 17224 26240
rect 17083 26200 17224 26228
rect 17083 26197 17095 26200
rect 17037 26191 17095 26197
rect 17218 26188 17224 26200
rect 17276 26188 17282 26240
rect 17402 26188 17408 26240
rect 17460 26228 17466 26240
rect 17880 26228 17908 26259
rect 20806 26256 20812 26268
rect 20864 26256 20870 26308
rect 18782 26228 18788 26240
rect 17460 26200 18788 26228
rect 17460 26188 17466 26200
rect 18782 26188 18788 26200
rect 18840 26188 18846 26240
rect 1104 26138 26312 26160
rect 1104 26086 4761 26138
rect 4813 26086 4825 26138
rect 4877 26086 4889 26138
rect 4941 26086 4953 26138
rect 5005 26086 5017 26138
rect 5069 26086 11063 26138
rect 11115 26086 11127 26138
rect 11179 26086 11191 26138
rect 11243 26086 11255 26138
rect 11307 26086 11319 26138
rect 11371 26086 17365 26138
rect 17417 26086 17429 26138
rect 17481 26086 17493 26138
rect 17545 26086 17557 26138
rect 17609 26086 17621 26138
rect 17673 26086 23667 26138
rect 23719 26086 23731 26138
rect 23783 26086 23795 26138
rect 23847 26086 23859 26138
rect 23911 26086 23923 26138
rect 23975 26086 26312 26138
rect 1104 26064 26312 26086
rect 9677 26027 9735 26033
rect 9677 26024 9689 26027
rect 6656 25996 9689 26024
rect 6546 25956 6552 25968
rect 6380 25928 6552 25956
rect 6380 25897 6408 25928
rect 6546 25916 6552 25928
rect 6604 25916 6610 25968
rect 6656 25965 6684 25996
rect 9677 25993 9689 25996
rect 9723 25993 9735 26027
rect 12802 26024 12808 26036
rect 9677 25987 9735 25993
rect 11532 25996 12808 26024
rect 6641 25959 6699 25965
rect 6641 25925 6653 25959
rect 6687 25925 6699 25959
rect 6641 25919 6699 25925
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 6972 25928 7130 25956
rect 6972 25916 6978 25928
rect 8938 25916 8944 25968
rect 8996 25956 9002 25968
rect 9309 25959 9367 25965
rect 8996 25928 9260 25956
rect 8996 25916 9002 25928
rect 6365 25891 6423 25897
rect 6365 25857 6377 25891
rect 6411 25857 6423 25891
rect 6365 25851 6423 25857
rect 8665 25891 8723 25897
rect 8665 25857 8677 25891
rect 8711 25857 8723 25891
rect 8665 25851 8723 25857
rect 8389 25823 8447 25829
rect 8389 25789 8401 25823
rect 8435 25820 8447 25823
rect 8680 25820 8708 25851
rect 9122 25848 9128 25900
rect 9180 25848 9186 25900
rect 9232 25888 9260 25928
rect 9309 25925 9321 25959
rect 9355 25956 9367 25959
rect 9582 25956 9588 25968
rect 9355 25928 9588 25956
rect 9355 25925 9367 25928
rect 9309 25919 9367 25925
rect 9582 25916 9588 25928
rect 9640 25916 9646 25968
rect 9876 25928 10548 25956
rect 9401 25891 9459 25897
rect 9401 25888 9413 25891
rect 9232 25860 9413 25888
rect 9401 25857 9413 25860
rect 9447 25857 9459 25891
rect 9401 25851 9459 25857
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25888 9551 25891
rect 9876 25888 9904 25928
rect 9539 25860 9904 25888
rect 9953 25891 10011 25897
rect 9539 25857 9551 25860
rect 9493 25851 9551 25857
rect 9953 25857 9965 25891
rect 9999 25857 10011 25891
rect 9953 25851 10011 25857
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 8435 25792 8708 25820
rect 8435 25789 8447 25792
rect 8389 25783 8447 25789
rect 8680 25752 8708 25792
rect 8754 25780 8760 25832
rect 8812 25780 8818 25832
rect 9033 25823 9091 25829
rect 9033 25789 9045 25823
rect 9079 25820 9091 25823
rect 9214 25820 9220 25832
rect 9079 25792 9220 25820
rect 9079 25789 9091 25792
rect 9033 25783 9091 25789
rect 9214 25780 9220 25792
rect 9272 25780 9278 25832
rect 9582 25780 9588 25832
rect 9640 25820 9646 25832
rect 9861 25823 9919 25829
rect 9861 25820 9873 25823
rect 9640 25792 9873 25820
rect 9640 25780 9646 25792
rect 9861 25789 9873 25792
rect 9907 25789 9919 25823
rect 9861 25783 9919 25789
rect 9968 25752 9996 25851
rect 10428 25820 10456 25851
rect 8680 25724 9996 25752
rect 10152 25792 10456 25820
rect 9232 25696 9260 25724
rect 9214 25644 9220 25696
rect 9272 25644 9278 25696
rect 9398 25644 9404 25696
rect 9456 25684 9462 25696
rect 10152 25684 10180 25792
rect 10321 25755 10379 25761
rect 10321 25721 10333 25755
rect 10367 25752 10379 25755
rect 10520 25752 10548 25928
rect 10594 25848 10600 25900
rect 10652 25848 10658 25900
rect 11532 25897 11560 25996
rect 12802 25984 12808 25996
rect 12860 25984 12866 26036
rect 13814 25984 13820 26036
rect 13872 25984 13878 26036
rect 14642 25984 14648 26036
rect 14700 26024 14706 26036
rect 15930 26024 15936 26036
rect 14700 25996 15936 26024
rect 14700 25984 14706 25996
rect 15930 25984 15936 25996
rect 15988 26024 15994 26036
rect 18690 26024 18696 26036
rect 15988 25996 18696 26024
rect 15988 25984 15994 25996
rect 12710 25916 12716 25968
rect 12768 25916 12774 25968
rect 15470 25916 15476 25968
rect 15528 25916 15534 25968
rect 11517 25891 11575 25897
rect 11517 25857 11529 25891
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 11793 25891 11851 25897
rect 11793 25857 11805 25891
rect 11839 25888 11851 25891
rect 11882 25888 11888 25900
rect 11839 25860 11888 25888
rect 11839 25857 11851 25860
rect 11793 25851 11851 25857
rect 11882 25848 11888 25860
rect 11940 25888 11946 25900
rect 11940 25860 12296 25888
rect 11940 25848 11946 25860
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 10367 25724 10548 25752
rect 11808 25792 12173 25820
rect 10367 25721 10379 25724
rect 10321 25715 10379 25721
rect 9456 25656 10180 25684
rect 9456 25644 9462 25656
rect 10226 25644 10232 25696
rect 10284 25684 10290 25696
rect 10413 25687 10471 25693
rect 10413 25684 10425 25687
rect 10284 25656 10425 25684
rect 10284 25644 10290 25656
rect 10413 25653 10425 25656
rect 10459 25653 10471 25687
rect 10413 25647 10471 25653
rect 11606 25644 11612 25696
rect 11664 25644 11670 25696
rect 11808 25684 11836 25792
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12268 25820 12296 25860
rect 13722 25848 13728 25900
rect 13780 25848 13786 25900
rect 16298 25848 16304 25900
rect 16356 25848 16362 25900
rect 16776 25897 16804 25996
rect 18690 25984 18696 25996
rect 18748 25984 18754 26036
rect 21913 26027 21971 26033
rect 21913 25993 21925 26027
rect 21959 26024 21971 26027
rect 23382 26024 23388 26036
rect 21959 25996 23388 26024
rect 21959 25993 21971 25996
rect 21913 25987 21971 25993
rect 23382 25984 23388 25996
rect 23440 25984 23446 26036
rect 19061 25959 19119 25965
rect 19061 25956 19073 25959
rect 18446 25928 19073 25956
rect 19061 25925 19073 25928
rect 19107 25925 19119 25959
rect 19061 25919 19119 25925
rect 20806 25916 20812 25968
rect 20864 25916 20870 25968
rect 23566 25916 23572 25968
rect 23624 25916 23630 25968
rect 16761 25891 16819 25897
rect 16761 25857 16773 25891
rect 16807 25857 16819 25891
rect 16761 25851 16819 25857
rect 17126 25848 17132 25900
rect 17184 25888 17190 25900
rect 17405 25891 17463 25897
rect 17405 25888 17417 25891
rect 17184 25860 17417 25888
rect 17184 25848 17190 25860
rect 17405 25857 17417 25860
rect 17451 25857 17463 25891
rect 17405 25851 17463 25857
rect 18969 25891 19027 25897
rect 18969 25857 18981 25891
rect 19015 25888 19027 25891
rect 19015 25860 19104 25888
rect 19015 25857 19027 25860
rect 18969 25851 19027 25857
rect 19076 25832 19104 25860
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19705 25891 19763 25897
rect 19705 25888 19717 25891
rect 19484 25860 19717 25888
rect 19484 25848 19490 25860
rect 19705 25857 19717 25860
rect 19751 25888 19763 25891
rect 19751 25860 20208 25888
rect 19751 25857 19763 25860
rect 19705 25851 19763 25857
rect 14369 25823 14427 25829
rect 14369 25820 14381 25823
rect 12268 25792 14381 25820
rect 12161 25783 12219 25789
rect 14369 25789 14381 25792
rect 14415 25789 14427 25823
rect 14369 25783 14427 25789
rect 14737 25823 14795 25829
rect 14737 25789 14749 25823
rect 14783 25820 14795 25823
rect 15470 25820 15476 25832
rect 14783 25792 15476 25820
rect 14783 25789 14795 25792
rect 14737 25783 14795 25789
rect 15470 25780 15476 25792
rect 15528 25780 15534 25832
rect 17034 25780 17040 25832
rect 17092 25780 17098 25832
rect 19058 25780 19064 25832
rect 19116 25780 19122 25832
rect 20070 25780 20076 25832
rect 20128 25780 20134 25832
rect 20180 25820 20208 25860
rect 22094 25848 22100 25900
rect 22152 25848 22158 25900
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25888 22247 25891
rect 22646 25888 22652 25900
rect 22235 25860 22652 25888
rect 22235 25857 22247 25860
rect 22189 25851 22247 25857
rect 22204 25820 22232 25851
rect 22646 25848 22652 25860
rect 22704 25848 22710 25900
rect 20180 25792 22232 25820
rect 22554 25780 22560 25832
rect 22612 25780 22618 25832
rect 15838 25712 15844 25764
rect 15896 25752 15902 25764
rect 16393 25755 16451 25761
rect 16393 25752 16405 25755
rect 15896 25724 16405 25752
rect 15896 25712 15902 25724
rect 16393 25721 16405 25724
rect 16439 25721 16451 25755
rect 16393 25715 16451 25721
rect 13446 25684 13452 25696
rect 11808 25656 13452 25684
rect 13446 25644 13452 25656
rect 13504 25644 13510 25696
rect 13541 25687 13599 25693
rect 13541 25653 13553 25687
rect 13587 25684 13599 25687
rect 13998 25684 14004 25696
rect 13587 25656 14004 25684
rect 13587 25653 13599 25656
rect 13541 25647 13599 25653
rect 13998 25644 14004 25656
rect 14056 25644 14062 25696
rect 16163 25687 16221 25693
rect 16163 25653 16175 25687
rect 16209 25684 16221 25687
rect 16298 25684 16304 25696
rect 16209 25656 16304 25684
rect 16209 25653 16221 25656
rect 16163 25647 16221 25653
rect 16298 25644 16304 25656
rect 16356 25644 16362 25696
rect 16853 25687 16911 25693
rect 16853 25653 16865 25687
rect 16899 25684 16911 25687
rect 18230 25684 18236 25696
rect 16899 25656 18236 25684
rect 16899 25653 16911 25656
rect 16853 25647 16911 25653
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 18782 25644 18788 25696
rect 18840 25644 18846 25696
rect 21266 25644 21272 25696
rect 21324 25684 21330 25696
rect 21453 25687 21511 25693
rect 21453 25684 21465 25687
rect 21324 25656 21465 25684
rect 21324 25644 21330 25656
rect 21453 25653 21465 25656
rect 21499 25653 21511 25687
rect 21453 25647 21511 25653
rect 23983 25687 24041 25693
rect 23983 25653 23995 25687
rect 24029 25684 24041 25687
rect 24394 25684 24400 25696
rect 24029 25656 24400 25684
rect 24029 25653 24041 25656
rect 23983 25647 24041 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 1104 25594 26312 25616
rect 1104 25542 4101 25594
rect 4153 25542 4165 25594
rect 4217 25542 4229 25594
rect 4281 25542 4293 25594
rect 4345 25542 4357 25594
rect 4409 25542 10403 25594
rect 10455 25542 10467 25594
rect 10519 25542 10531 25594
rect 10583 25542 10595 25594
rect 10647 25542 10659 25594
rect 10711 25542 16705 25594
rect 16757 25542 16769 25594
rect 16821 25542 16833 25594
rect 16885 25542 16897 25594
rect 16949 25542 16961 25594
rect 17013 25542 23007 25594
rect 23059 25542 23071 25594
rect 23123 25542 23135 25594
rect 23187 25542 23199 25594
rect 23251 25542 23263 25594
rect 23315 25542 26312 25594
rect 1104 25520 26312 25542
rect 6914 25440 6920 25492
rect 6972 25440 6978 25492
rect 7466 25440 7472 25492
rect 7524 25440 7530 25492
rect 9030 25440 9036 25492
rect 9088 25480 9094 25492
rect 9769 25483 9827 25489
rect 9088 25452 9674 25480
rect 9088 25440 9094 25452
rect 9125 25415 9183 25421
rect 9125 25381 9137 25415
rect 9171 25412 9183 25415
rect 9646 25412 9674 25452
rect 9769 25449 9781 25483
rect 9815 25480 9827 25483
rect 9950 25480 9956 25492
rect 9815 25452 9956 25480
rect 9815 25449 9827 25452
rect 9769 25443 9827 25449
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 12710 25440 12716 25492
rect 12768 25440 12774 25492
rect 12802 25440 12808 25492
rect 12860 25480 12866 25492
rect 13722 25480 13728 25492
rect 12860 25452 13728 25480
rect 12860 25440 12866 25452
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 15470 25440 15476 25492
rect 15528 25440 15534 25492
rect 17862 25480 17868 25492
rect 16960 25452 17868 25480
rect 9171 25384 9536 25412
rect 9646 25384 9812 25412
rect 9171 25381 9183 25384
rect 9125 25375 9183 25381
rect 4709 25347 4767 25353
rect 4709 25313 4721 25347
rect 4755 25344 4767 25347
rect 6546 25344 6552 25356
rect 4755 25316 6552 25344
rect 4755 25313 4767 25316
rect 4709 25307 4767 25313
rect 6546 25304 6552 25316
rect 6604 25304 6610 25356
rect 8294 25304 8300 25356
rect 8352 25344 8358 25356
rect 9508 25344 9536 25384
rect 9784 25356 9812 25384
rect 9858 25372 9864 25424
rect 9916 25372 9922 25424
rect 10226 25372 10232 25424
rect 10284 25372 10290 25424
rect 12434 25372 12440 25424
rect 12492 25412 12498 25424
rect 13078 25412 13084 25424
rect 12492 25384 13084 25412
rect 12492 25372 12498 25384
rect 13078 25372 13084 25384
rect 13136 25412 13142 25424
rect 13265 25415 13323 25421
rect 13265 25412 13277 25415
rect 13136 25384 13277 25412
rect 13136 25372 13142 25384
rect 13265 25381 13277 25384
rect 13311 25381 13323 25415
rect 13265 25375 13323 25381
rect 13538 25372 13544 25424
rect 13596 25372 13602 25424
rect 14844 25384 15792 25412
rect 8352 25316 9352 25344
rect 9508 25316 9628 25344
rect 8352 25304 8358 25316
rect 6822 25236 6828 25288
rect 6880 25276 6886 25288
rect 7377 25279 7435 25285
rect 7377 25276 7389 25279
rect 6880 25248 7389 25276
rect 6880 25236 6886 25248
rect 7377 25245 7389 25248
rect 7423 25245 7435 25279
rect 7377 25239 7435 25245
rect 9122 25236 9128 25288
rect 9180 25236 9186 25288
rect 9324 25285 9352 25316
rect 9600 25288 9628 25316
rect 9766 25304 9772 25356
rect 9824 25304 9830 25356
rect 10244 25344 10272 25372
rect 14844 25356 14872 25384
rect 10505 25347 10563 25353
rect 10505 25344 10517 25347
rect 10060 25316 10517 25344
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25276 9367 25279
rect 9490 25276 9496 25288
rect 9355 25248 9496 25276
rect 9355 25245 9367 25248
rect 9309 25239 9367 25245
rect 9490 25236 9496 25248
rect 9548 25236 9554 25288
rect 9582 25236 9588 25288
rect 9640 25236 9646 25288
rect 9674 25236 9680 25288
rect 9732 25276 9738 25288
rect 10060 25285 10088 25316
rect 10505 25313 10517 25316
rect 10551 25313 10563 25347
rect 10505 25307 10563 25313
rect 10870 25304 10876 25356
rect 10928 25344 10934 25356
rect 12253 25347 12311 25353
rect 12253 25344 12265 25347
rect 10928 25316 12265 25344
rect 10928 25304 10934 25316
rect 12253 25313 12265 25316
rect 12299 25313 12311 25347
rect 14826 25344 14832 25356
rect 12253 25307 12311 25313
rect 13280 25316 14832 25344
rect 9861 25279 9919 25285
rect 9861 25276 9873 25279
rect 9732 25248 9873 25276
rect 9732 25236 9738 25248
rect 9861 25245 9873 25248
rect 9907 25245 9919 25279
rect 9861 25239 9919 25245
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25245 10103 25279
rect 10045 25239 10103 25245
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 4985 25211 5043 25217
rect 4985 25177 4997 25211
rect 5031 25177 5043 25211
rect 4985 25171 5043 25177
rect 5000 25140 5028 25171
rect 5994 25168 6000 25220
rect 6052 25168 6058 25220
rect 6730 25168 6736 25220
rect 6788 25168 6794 25220
rect 8754 25168 8760 25220
rect 8812 25208 8818 25220
rect 9398 25208 9404 25220
rect 8812 25180 9404 25208
rect 8812 25168 8818 25180
rect 9398 25168 9404 25180
rect 9456 25168 9462 25220
rect 9950 25168 9956 25220
rect 10008 25208 10014 25220
rect 10152 25208 10180 25239
rect 10226 25236 10232 25288
rect 10284 25236 10290 25288
rect 11606 25236 11612 25288
rect 11664 25236 11670 25288
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25276 12679 25279
rect 12802 25276 12808 25288
rect 12667 25248 12808 25276
rect 12667 25245 12679 25248
rect 12621 25239 12679 25245
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 13280 25285 13308 25316
rect 14826 25304 14832 25316
rect 14884 25304 14890 25356
rect 15565 25347 15623 25353
rect 15565 25344 15577 25347
rect 15120 25316 15577 25344
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25245 13323 25279
rect 13265 25239 13323 25245
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25245 13507 25279
rect 13449 25239 13507 25245
rect 10008 25180 10180 25208
rect 10008 25168 10014 25180
rect 6454 25140 6460 25152
rect 5000 25112 6460 25140
rect 6454 25100 6460 25112
rect 6512 25100 6518 25152
rect 6546 25100 6552 25152
rect 6604 25140 6610 25152
rect 10226 25140 10232 25152
rect 6604 25112 10232 25140
rect 6604 25100 6610 25112
rect 10226 25100 10232 25112
rect 10284 25100 10290 25152
rect 13464 25140 13492 25239
rect 13814 25236 13820 25288
rect 13872 25236 13878 25288
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25276 14611 25279
rect 14642 25276 14648 25288
rect 14599 25248 14648 25276
rect 14599 25245 14611 25248
rect 14553 25239 14611 25245
rect 14642 25236 14648 25248
rect 14700 25236 14706 25288
rect 14918 25236 14924 25288
rect 14976 25236 14982 25288
rect 15120 25285 15148 25316
rect 15565 25313 15577 25316
rect 15611 25313 15623 25347
rect 15565 25307 15623 25313
rect 15764 25288 15792 25384
rect 16390 25304 16396 25356
rect 16448 25344 16454 25356
rect 16761 25347 16819 25353
rect 16761 25344 16773 25347
rect 16448 25316 16773 25344
rect 16448 25304 16454 25316
rect 16761 25313 16773 25316
rect 16807 25344 16819 25347
rect 16960 25344 16988 25452
rect 17862 25440 17868 25452
rect 17920 25440 17926 25492
rect 23566 25440 23572 25492
rect 23624 25480 23630 25492
rect 23661 25483 23719 25489
rect 23661 25480 23673 25483
rect 23624 25452 23673 25480
rect 23624 25440 23630 25452
rect 23661 25449 23673 25452
rect 23707 25449 23719 25483
rect 23661 25443 23719 25449
rect 20806 25372 20812 25424
rect 20864 25412 20870 25424
rect 23017 25415 23075 25421
rect 23017 25412 23029 25415
rect 20864 25384 23029 25412
rect 20864 25372 20870 25384
rect 23017 25381 23029 25384
rect 23063 25381 23075 25415
rect 23017 25375 23075 25381
rect 16807 25316 16988 25344
rect 16807 25313 16819 25316
rect 16761 25307 16819 25313
rect 17034 25304 17040 25356
rect 17092 25344 17098 25356
rect 17129 25347 17187 25353
rect 17129 25344 17141 25347
rect 17092 25316 17141 25344
rect 17092 25304 17098 25316
rect 17129 25313 17141 25316
rect 17175 25344 17187 25347
rect 19426 25344 19432 25356
rect 17175 25316 19432 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 19426 25304 19432 25316
rect 19484 25304 19490 25356
rect 21358 25304 21364 25356
rect 21416 25304 21422 25356
rect 22066 25316 23336 25344
rect 22066 25288 22094 25316
rect 15105 25279 15163 25285
rect 15105 25245 15117 25279
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 15286 25236 15292 25288
rect 15344 25236 15350 25288
rect 15746 25236 15752 25288
rect 15804 25236 15810 25288
rect 16022 25236 16028 25288
rect 16080 25236 16086 25288
rect 16669 25279 16727 25285
rect 16669 25245 16681 25279
rect 16715 25276 16727 25279
rect 16942 25276 16948 25288
rect 16715 25248 16948 25276
rect 16715 25245 16727 25248
rect 16669 25239 16727 25245
rect 16942 25236 16948 25248
rect 17000 25236 17006 25288
rect 17218 25236 17224 25288
rect 17276 25276 17282 25288
rect 17497 25279 17555 25285
rect 17497 25276 17509 25279
rect 17276 25248 17509 25276
rect 17276 25236 17282 25248
rect 17497 25245 17509 25248
rect 17543 25245 17555 25279
rect 17497 25239 17555 25245
rect 21266 25236 21272 25288
rect 21324 25276 21330 25288
rect 21453 25279 21511 25285
rect 21453 25276 21465 25279
rect 21324 25248 21465 25276
rect 21324 25236 21330 25248
rect 21453 25245 21465 25248
rect 21499 25276 21511 25279
rect 22002 25276 22008 25288
rect 21499 25248 22008 25276
rect 21499 25245 21511 25248
rect 21453 25239 21511 25245
rect 22002 25236 22008 25248
rect 22060 25248 22094 25288
rect 22060 25236 22066 25248
rect 22462 25236 22468 25288
rect 22520 25276 22526 25288
rect 23308 25285 23336 25316
rect 23293 25279 23351 25285
rect 22520 25248 23244 25276
rect 22520 25236 22526 25248
rect 13541 25211 13599 25217
rect 13541 25177 13553 25211
rect 13587 25208 13599 25211
rect 13587 25180 14780 25208
rect 13587 25177 13599 25180
rect 13541 25171 13599 25177
rect 13725 25143 13783 25149
rect 13725 25140 13737 25143
rect 13464 25112 13737 25140
rect 13725 25109 13737 25112
rect 13771 25140 13783 25143
rect 14366 25140 14372 25152
rect 13771 25112 14372 25140
rect 13771 25109 13783 25112
rect 13725 25103 13783 25109
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 14752 25149 14780 25180
rect 15010 25168 15016 25220
rect 15068 25208 15074 25220
rect 15197 25211 15255 25217
rect 15197 25208 15209 25211
rect 15068 25180 15209 25208
rect 15068 25168 15074 25180
rect 15197 25177 15209 25180
rect 15243 25208 15255 25211
rect 19150 25208 19156 25220
rect 15243 25180 17264 25208
rect 18538 25180 19156 25208
rect 15243 25177 15255 25180
rect 15197 25171 15255 25177
rect 17236 25152 17264 25180
rect 19150 25168 19156 25180
rect 19208 25168 19214 25220
rect 19702 25168 19708 25220
rect 19760 25168 19766 25220
rect 20714 25168 20720 25220
rect 20772 25168 20778 25220
rect 21358 25168 21364 25220
rect 21416 25208 21422 25220
rect 23109 25211 23167 25217
rect 23109 25208 23121 25211
rect 21416 25180 23121 25208
rect 21416 25168 21422 25180
rect 23109 25177 23121 25180
rect 23155 25177 23167 25211
rect 23216 25208 23244 25248
rect 23293 25245 23305 25279
rect 23339 25245 23351 25279
rect 23293 25239 23351 25245
rect 23569 25279 23627 25285
rect 23569 25245 23581 25279
rect 23615 25276 23627 25279
rect 24302 25276 24308 25288
rect 23615 25248 24308 25276
rect 23615 25245 23627 25248
rect 23569 25239 23627 25245
rect 24302 25236 24308 25248
rect 24360 25236 24366 25288
rect 24394 25236 24400 25288
rect 24452 25236 24458 25288
rect 25774 25236 25780 25288
rect 25832 25236 25838 25288
rect 24412 25208 24440 25236
rect 23216 25180 24440 25208
rect 23109 25171 23167 25177
rect 14737 25143 14795 25149
rect 14737 25109 14749 25143
rect 14783 25140 14795 25143
rect 14918 25140 14924 25152
rect 14783 25112 14924 25140
rect 14783 25109 14795 25112
rect 14737 25103 14795 25109
rect 14918 25100 14924 25112
rect 14976 25100 14982 25152
rect 15933 25143 15991 25149
rect 15933 25109 15945 25143
rect 15979 25140 15991 25143
rect 16758 25140 16764 25152
rect 15979 25112 16764 25140
rect 15979 25109 15991 25112
rect 15933 25103 15991 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 17034 25100 17040 25152
rect 17092 25100 17098 25152
rect 17218 25100 17224 25152
rect 17276 25100 17282 25152
rect 18874 25100 18880 25152
rect 18932 25149 18938 25152
rect 18932 25143 18981 25149
rect 18932 25109 18935 25143
rect 18969 25109 18981 25143
rect 18932 25103 18981 25109
rect 18932 25100 18938 25103
rect 21174 25100 21180 25152
rect 21232 25100 21238 25152
rect 21818 25100 21824 25152
rect 21876 25100 21882 25152
rect 22094 25100 22100 25152
rect 22152 25140 22158 25152
rect 22738 25140 22744 25152
rect 22152 25112 22744 25140
rect 22152 25100 22158 25112
rect 22738 25100 22744 25112
rect 22796 25100 22802 25152
rect 23474 25100 23480 25152
rect 23532 25100 23538 25152
rect 25038 25100 25044 25152
rect 25096 25100 25102 25152
rect 25222 25100 25228 25152
rect 25280 25140 25286 25152
rect 25961 25143 26019 25149
rect 25961 25140 25973 25143
rect 25280 25112 25973 25140
rect 25280 25100 25286 25112
rect 25961 25109 25973 25112
rect 26007 25109 26019 25143
rect 25961 25103 26019 25109
rect 1104 25050 26312 25072
rect 1104 24998 4761 25050
rect 4813 24998 4825 25050
rect 4877 24998 4889 25050
rect 4941 24998 4953 25050
rect 5005 24998 5017 25050
rect 5069 24998 11063 25050
rect 11115 24998 11127 25050
rect 11179 24998 11191 25050
rect 11243 24998 11255 25050
rect 11307 24998 11319 25050
rect 11371 24998 17365 25050
rect 17417 24998 17429 25050
rect 17481 24998 17493 25050
rect 17545 24998 17557 25050
rect 17609 24998 17621 25050
rect 17673 24998 23667 25050
rect 23719 24998 23731 25050
rect 23783 24998 23795 25050
rect 23847 24998 23859 25050
rect 23911 24998 23923 25050
rect 23975 24998 26312 25050
rect 1104 24976 26312 24998
rect 7101 24939 7159 24945
rect 7101 24905 7113 24939
rect 7147 24936 7159 24939
rect 8110 24936 8116 24948
rect 7147 24908 8116 24936
rect 7147 24905 7159 24908
rect 7101 24899 7159 24905
rect 8110 24896 8116 24908
rect 8168 24896 8174 24948
rect 9398 24896 9404 24948
rect 9456 24945 9462 24948
rect 9456 24939 9475 24945
rect 9463 24936 9475 24939
rect 9463 24908 9536 24936
rect 9463 24905 9475 24908
rect 9456 24899 9475 24905
rect 9456 24896 9462 24899
rect 6822 24868 6828 24880
rect 5828 24840 6828 24868
rect 5828 24809 5856 24840
rect 6822 24828 6828 24840
rect 6880 24828 6886 24880
rect 9217 24871 9275 24877
rect 7300 24840 7512 24868
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24769 5871 24803
rect 5813 24763 5871 24769
rect 5905 24803 5963 24809
rect 5905 24769 5917 24803
rect 5951 24800 5963 24803
rect 5994 24800 6000 24812
rect 5951 24772 6000 24800
rect 5951 24769 5963 24772
rect 5905 24763 5963 24769
rect 5994 24760 6000 24772
rect 6052 24760 6058 24812
rect 6730 24760 6736 24812
rect 6788 24760 6794 24812
rect 7300 24800 7328 24840
rect 6840 24772 7328 24800
rect 7377 24803 7435 24809
rect 6748 24664 6776 24760
rect 6840 24741 6868 24772
rect 7377 24769 7389 24803
rect 7423 24769 7435 24803
rect 7484 24800 7512 24840
rect 7760 24840 8984 24868
rect 7558 24800 7564 24812
rect 7484 24772 7564 24800
rect 7377 24763 7435 24769
rect 6825 24735 6883 24741
rect 6825 24701 6837 24735
rect 6871 24701 6883 24735
rect 6825 24695 6883 24701
rect 7392 24664 7420 24763
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 7650 24760 7656 24812
rect 7708 24760 7714 24812
rect 7760 24732 7788 24840
rect 7834 24760 7840 24812
rect 7892 24760 7898 24812
rect 8018 24760 8024 24812
rect 8076 24760 8082 24812
rect 8956 24809 8984 24840
rect 9217 24837 9229 24871
rect 9263 24837 9275 24871
rect 9217 24831 9275 24837
rect 8389 24803 8447 24809
rect 8389 24769 8401 24803
rect 8435 24769 8447 24803
rect 8389 24763 8447 24769
rect 8941 24803 8999 24809
rect 8941 24769 8953 24803
rect 8987 24800 8999 24803
rect 9030 24800 9036 24812
rect 8987 24772 9036 24800
rect 8987 24769 8999 24772
rect 8941 24763 8999 24769
rect 7484 24704 7788 24732
rect 7852 24732 7880 24760
rect 8294 24732 8300 24744
rect 7852 24704 8300 24732
rect 7484 24676 7512 24704
rect 8294 24692 8300 24704
rect 8352 24732 8358 24744
rect 8404 24732 8432 24763
rect 9030 24760 9036 24772
rect 9088 24760 9094 24812
rect 8352 24704 8432 24732
rect 9232 24732 9260 24831
rect 9508 24800 9536 24908
rect 13078 24896 13084 24948
rect 13136 24896 13142 24948
rect 13814 24896 13820 24948
rect 13872 24936 13878 24948
rect 14001 24939 14059 24945
rect 14001 24936 14013 24939
rect 13872 24908 14013 24936
rect 13872 24896 13878 24908
rect 14001 24905 14013 24908
rect 14047 24905 14059 24939
rect 14918 24936 14924 24948
rect 14001 24899 14059 24905
rect 14108 24908 14924 24936
rect 12897 24871 12955 24877
rect 12897 24837 12909 24871
rect 12943 24868 12955 24871
rect 13538 24868 13544 24880
rect 12943 24840 13544 24868
rect 12943 24837 12955 24840
rect 12897 24831 12955 24837
rect 13538 24828 13544 24840
rect 13596 24828 13602 24880
rect 13832 24868 13860 24896
rect 13740 24840 13860 24868
rect 9861 24803 9919 24809
rect 9508 24772 9812 24800
rect 9232 24704 9628 24732
rect 8352 24692 8358 24704
rect 6748 24636 7420 24664
rect 7193 24599 7251 24605
rect 7193 24565 7205 24599
rect 7239 24596 7251 24599
rect 7282 24596 7288 24608
rect 7239 24568 7288 24596
rect 7239 24565 7251 24568
rect 7193 24559 7251 24565
rect 7282 24556 7288 24568
rect 7340 24556 7346 24608
rect 7392 24596 7420 24636
rect 7466 24624 7472 24676
rect 7524 24624 7530 24676
rect 8018 24664 8024 24676
rect 7576 24636 8024 24664
rect 7576 24596 7604 24636
rect 8018 24624 8024 24636
rect 8076 24624 8082 24676
rect 8404 24664 8432 24704
rect 9600 24664 9628 24704
rect 9674 24692 9680 24744
rect 9732 24692 9738 24744
rect 9784 24732 9812 24772
rect 9861 24769 9873 24803
rect 9907 24800 9919 24803
rect 10134 24800 10140 24812
rect 9907 24772 10140 24800
rect 9907 24769 9919 24772
rect 9861 24763 9919 24769
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 13173 24803 13231 24809
rect 13173 24769 13185 24803
rect 13219 24769 13231 24803
rect 13173 24763 13231 24769
rect 10045 24735 10103 24741
rect 10045 24732 10057 24735
rect 9784 24704 10057 24732
rect 10045 24701 10057 24704
rect 10091 24701 10103 24735
rect 13188 24732 13216 24763
rect 13630 24760 13636 24812
rect 13688 24760 13694 24812
rect 13740 24732 13768 24840
rect 13817 24803 13875 24809
rect 13817 24769 13829 24803
rect 13863 24800 13875 24803
rect 13906 24800 13912 24812
rect 13863 24772 13912 24800
rect 13863 24769 13875 24772
rect 13817 24763 13875 24769
rect 13906 24760 13912 24772
rect 13964 24760 13970 24812
rect 14108 24809 14136 24908
rect 14918 24896 14924 24908
rect 14976 24896 14982 24948
rect 15286 24896 15292 24948
rect 15344 24936 15350 24948
rect 15473 24939 15531 24945
rect 15473 24936 15485 24939
rect 15344 24908 15485 24936
rect 15344 24896 15350 24908
rect 15473 24905 15485 24908
rect 15519 24905 15531 24939
rect 15473 24899 15531 24905
rect 15746 24896 15752 24948
rect 15804 24936 15810 24948
rect 16485 24939 16543 24945
rect 16485 24936 16497 24939
rect 15804 24908 16497 24936
rect 15804 24896 15810 24908
rect 16485 24905 16497 24908
rect 16531 24905 16543 24939
rect 16485 24899 16543 24905
rect 16574 24896 16580 24948
rect 16632 24896 16638 24948
rect 16945 24939 17003 24945
rect 16945 24905 16957 24939
rect 16991 24936 17003 24939
rect 17126 24936 17132 24948
rect 16991 24908 17132 24936
rect 16991 24905 17003 24908
rect 16945 24899 17003 24905
rect 17126 24896 17132 24908
rect 17184 24896 17190 24948
rect 17218 24896 17224 24948
rect 17276 24936 17282 24948
rect 17773 24939 17831 24945
rect 17773 24936 17785 24939
rect 17276 24908 17785 24936
rect 17276 24896 17282 24908
rect 14366 24828 14372 24880
rect 14424 24868 14430 24880
rect 15010 24868 15016 24880
rect 14424 24840 15016 24868
rect 14424 24828 14430 24840
rect 15010 24828 15016 24840
rect 15068 24828 15074 24880
rect 16117 24871 16175 24877
rect 16117 24837 16129 24871
rect 16163 24868 16175 24871
rect 16333 24871 16391 24877
rect 16163 24840 16252 24868
rect 16163 24837 16175 24840
rect 16117 24831 16175 24837
rect 14093 24803 14151 24809
rect 14093 24769 14105 24803
rect 14139 24769 14151 24803
rect 14093 24763 14151 24769
rect 14277 24803 14335 24809
rect 14277 24769 14289 24803
rect 14323 24769 14335 24803
rect 14277 24763 14335 24769
rect 13188 24704 13768 24732
rect 14292 24732 14320 24763
rect 14458 24760 14464 24812
rect 14516 24760 14522 24812
rect 14642 24760 14648 24812
rect 14700 24800 14706 24812
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 14700 24772 14749 24800
rect 14700 24760 14706 24772
rect 14737 24769 14749 24772
rect 14783 24769 14795 24803
rect 14737 24763 14795 24769
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 14921 24803 14979 24809
rect 14921 24800 14933 24803
rect 14884 24772 14933 24800
rect 14884 24760 14890 24772
rect 14921 24769 14933 24772
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15381 24803 15439 24809
rect 15381 24800 15393 24803
rect 15252 24772 15393 24800
rect 15252 24760 15258 24772
rect 15381 24769 15393 24772
rect 15427 24769 15439 24803
rect 15381 24763 15439 24769
rect 15565 24803 15623 24809
rect 15565 24769 15577 24803
rect 15611 24769 15623 24803
rect 16224 24800 16252 24840
rect 16333 24837 16345 24871
rect 16379 24868 16391 24871
rect 16592 24868 16620 24896
rect 17446 24877 17474 24908
rect 17773 24905 17785 24908
rect 17819 24905 17831 24939
rect 17773 24899 17831 24905
rect 19702 24896 19708 24948
rect 19760 24896 19766 24948
rect 20070 24896 20076 24948
rect 20128 24936 20134 24948
rect 20349 24939 20407 24945
rect 20349 24936 20361 24939
rect 20128 24908 20361 24936
rect 20128 24896 20134 24908
rect 20349 24905 20361 24908
rect 20395 24905 20407 24939
rect 22186 24936 22192 24948
rect 20349 24899 20407 24905
rect 20456 24908 22192 24936
rect 17431 24871 17489 24877
rect 16379 24840 16712 24868
rect 16379 24837 16391 24840
rect 16333 24831 16391 24837
rect 16574 24800 16580 24812
rect 16224 24772 16580 24800
rect 15565 24763 15623 24769
rect 15105 24735 15163 24741
rect 15105 24732 15117 24735
rect 14292 24704 15117 24732
rect 10045 24695 10103 24701
rect 15105 24701 15117 24704
rect 15151 24701 15163 24735
rect 15580 24732 15608 24763
rect 16574 24760 16580 24772
rect 16632 24760 16638 24812
rect 16684 24809 16712 24840
rect 17431 24837 17443 24871
rect 17477 24837 17489 24871
rect 18782 24868 18788 24880
rect 17431 24831 17489 24837
rect 18156 24840 18788 24868
rect 18156 24812 18184 24840
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 15746 24732 15752 24744
rect 15580 24704 15752 24732
rect 15105 24695 15163 24701
rect 15746 24692 15752 24704
rect 15804 24732 15810 24744
rect 16390 24732 16396 24744
rect 15804 24704 16396 24732
rect 15804 24692 15810 24704
rect 16390 24692 16396 24704
rect 16448 24692 16454 24744
rect 16482 24692 16488 24744
rect 16540 24732 16546 24744
rect 16684 24732 16712 24763
rect 16758 24760 16764 24812
rect 16816 24760 16822 24812
rect 17034 24760 17040 24812
rect 17092 24760 17098 24812
rect 17126 24760 17132 24812
rect 17184 24760 17190 24812
rect 17218 24760 17224 24812
rect 17276 24760 17282 24812
rect 17310 24760 17316 24812
rect 17368 24760 17374 24812
rect 17954 24760 17960 24812
rect 18012 24760 18018 24812
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24800 18107 24803
rect 18138 24800 18144 24812
rect 18095 24772 18144 24800
rect 18095 24769 18107 24772
rect 18049 24763 18107 24769
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 18230 24760 18236 24812
rect 18288 24760 18294 24812
rect 18414 24760 18420 24812
rect 18472 24760 18478 24812
rect 18616 24809 18644 24840
rect 18782 24828 18788 24840
rect 18840 24828 18846 24880
rect 18601 24803 18659 24809
rect 18601 24769 18613 24803
rect 18647 24769 18659 24803
rect 18601 24763 18659 24769
rect 18690 24760 18696 24812
rect 18748 24760 18754 24812
rect 18874 24760 18880 24812
rect 18932 24760 18938 24812
rect 19058 24760 19064 24812
rect 19116 24760 19122 24812
rect 19150 24760 19156 24812
rect 19208 24760 19214 24812
rect 19981 24803 20039 24809
rect 19981 24769 19993 24803
rect 20027 24800 20039 24803
rect 20456 24800 20484 24908
rect 22186 24896 22192 24908
rect 22244 24936 22250 24948
rect 22462 24936 22468 24948
rect 22244 24908 22468 24936
rect 22244 24896 22250 24908
rect 22462 24896 22468 24908
rect 22520 24896 22526 24948
rect 20714 24828 20720 24880
rect 20772 24828 20778 24880
rect 21818 24868 21824 24880
rect 21008 24840 21824 24868
rect 20027 24772 20484 24800
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 20530 24760 20536 24812
rect 20588 24760 20594 24812
rect 20622 24760 20628 24812
rect 20680 24760 20686 24812
rect 20806 24760 20812 24812
rect 20864 24809 20870 24812
rect 21008 24809 21036 24840
rect 21818 24828 21824 24840
rect 21876 24828 21882 24880
rect 20864 24803 20893 24809
rect 20881 24769 20893 24803
rect 20864 24763 20893 24769
rect 20993 24803 21051 24809
rect 20993 24769 21005 24803
rect 21039 24769 21051 24803
rect 20993 24763 21051 24769
rect 20864 24760 20870 24763
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 21269 24803 21327 24809
rect 21269 24800 21281 24803
rect 21232 24772 21281 24800
rect 21232 24760 21238 24772
rect 21269 24769 21281 24772
rect 21315 24769 21327 24803
rect 21269 24763 21327 24769
rect 21545 24803 21603 24809
rect 21545 24769 21557 24803
rect 21591 24769 21603 24803
rect 21545 24763 21603 24769
rect 16540 24704 16712 24732
rect 16540 24692 16546 24704
rect 10318 24664 10324 24676
rect 8404 24636 9536 24664
rect 9600 24636 10324 24664
rect 7392 24568 7604 24596
rect 8202 24556 8208 24608
rect 8260 24556 8266 24608
rect 8478 24556 8484 24608
rect 8536 24556 8542 24608
rect 8938 24556 8944 24608
rect 8996 24596 9002 24608
rect 9033 24599 9091 24605
rect 9033 24596 9045 24599
rect 8996 24568 9045 24596
rect 8996 24556 9002 24568
rect 9033 24565 9045 24568
rect 9079 24565 9091 24599
rect 9033 24559 9091 24565
rect 9214 24556 9220 24608
rect 9272 24596 9278 24608
rect 9401 24599 9459 24605
rect 9401 24596 9413 24599
rect 9272 24568 9413 24596
rect 9272 24556 9278 24568
rect 9401 24565 9413 24568
rect 9447 24565 9459 24599
rect 9508 24596 9536 24636
rect 9692 24608 9720 24636
rect 10318 24624 10324 24636
rect 10376 24624 10382 24676
rect 13446 24624 13452 24676
rect 13504 24664 13510 24676
rect 14645 24667 14703 24673
rect 14645 24664 14657 24667
rect 13504 24636 14657 24664
rect 13504 24624 13510 24636
rect 14645 24633 14657 24636
rect 14691 24633 14703 24667
rect 14645 24627 14703 24633
rect 14918 24624 14924 24676
rect 14976 24664 14982 24676
rect 16776 24664 16804 24760
rect 17052 24732 17080 24760
rect 17589 24735 17647 24741
rect 17589 24732 17601 24735
rect 17052 24704 17601 24732
rect 17589 24701 17601 24704
rect 17635 24701 17647 24735
rect 17972 24732 18000 24760
rect 18892 24732 18920 24760
rect 17972 24704 18920 24732
rect 17589 24695 17647 24701
rect 19886 24692 19892 24744
rect 19944 24692 19950 24744
rect 20070 24692 20076 24744
rect 20128 24692 20134 24744
rect 20165 24735 20223 24741
rect 20165 24701 20177 24735
rect 20211 24701 20223 24735
rect 21549 24732 21577 24763
rect 22094 24760 22100 24812
rect 22152 24760 22158 24812
rect 22186 24760 22192 24812
rect 22244 24760 22250 24812
rect 22370 24760 22376 24812
rect 22428 24760 22434 24812
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 22557 24803 22615 24809
rect 22557 24800 22569 24803
rect 22520 24772 22569 24800
rect 22520 24760 22526 24772
rect 22557 24769 22569 24772
rect 22603 24769 22615 24803
rect 22557 24763 22615 24769
rect 22649 24735 22707 24741
rect 22649 24732 22661 24735
rect 21549 24704 22661 24732
rect 20165 24695 20223 24701
rect 22649 24701 22661 24704
rect 22695 24701 22707 24735
rect 22649 24695 22707 24701
rect 17494 24664 17500 24676
rect 14976 24636 16620 24664
rect 16776 24636 17500 24664
rect 14976 24624 14982 24636
rect 9585 24599 9643 24605
rect 9585 24596 9597 24599
rect 9508 24568 9597 24596
rect 9401 24559 9459 24565
rect 9585 24565 9597 24568
rect 9631 24565 9643 24599
rect 9585 24559 9643 24565
rect 9674 24556 9680 24608
rect 9732 24556 9738 24608
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 12897 24599 12955 24605
rect 12897 24596 12909 24599
rect 12492 24568 12909 24596
rect 12492 24556 12498 24568
rect 12897 24565 12909 24568
rect 12943 24565 12955 24599
rect 12897 24559 12955 24565
rect 16301 24599 16359 24605
rect 16301 24565 16313 24599
rect 16347 24596 16359 24599
rect 16390 24596 16396 24608
rect 16347 24568 16396 24596
rect 16347 24565 16359 24568
rect 16301 24559 16359 24565
rect 16390 24556 16396 24568
rect 16448 24556 16454 24608
rect 16592 24596 16620 24636
rect 17494 24624 17500 24636
rect 17552 24624 17558 24676
rect 17862 24624 17868 24676
rect 17920 24664 17926 24676
rect 18141 24667 18199 24673
rect 18141 24664 18153 24667
rect 17920 24636 18153 24664
rect 17920 24624 17926 24636
rect 18141 24633 18153 24636
rect 18187 24633 18199 24667
rect 18141 24627 18199 24633
rect 18785 24667 18843 24673
rect 18785 24633 18797 24667
rect 18831 24633 18843 24667
rect 20180 24664 20208 24695
rect 20180 24636 21220 24664
rect 18785 24627 18843 24633
rect 17310 24596 17316 24608
rect 16592 24568 17316 24596
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 18156 24596 18184 24627
rect 18800 24596 18828 24627
rect 18156 24568 18828 24596
rect 20806 24556 20812 24608
rect 20864 24596 20870 24608
rect 21085 24599 21143 24605
rect 21085 24596 21097 24599
rect 20864 24568 21097 24596
rect 20864 24556 20870 24568
rect 21085 24565 21097 24568
rect 21131 24565 21143 24599
rect 21192 24596 21220 24636
rect 21266 24624 21272 24676
rect 21324 24664 21330 24676
rect 21361 24667 21419 24673
rect 21361 24664 21373 24667
rect 21324 24636 21373 24664
rect 21324 24624 21330 24636
rect 21361 24633 21373 24636
rect 21407 24633 21419 24667
rect 21361 24627 21419 24633
rect 21450 24624 21456 24676
rect 21508 24664 21514 24676
rect 22281 24667 22339 24673
rect 21508 24636 22094 24664
rect 21508 24624 21514 24636
rect 21913 24599 21971 24605
rect 21913 24596 21925 24599
rect 21192 24568 21925 24596
rect 21085 24559 21143 24565
rect 21913 24565 21925 24568
rect 21959 24565 21971 24599
rect 22066 24596 22094 24636
rect 22281 24633 22293 24667
rect 22327 24633 22339 24667
rect 22281 24627 22339 24633
rect 22296 24596 22324 24627
rect 22066 24568 22324 24596
rect 21913 24559 21971 24565
rect 1104 24506 26312 24528
rect 1104 24454 4101 24506
rect 4153 24454 4165 24506
rect 4217 24454 4229 24506
rect 4281 24454 4293 24506
rect 4345 24454 4357 24506
rect 4409 24454 10403 24506
rect 10455 24454 10467 24506
rect 10519 24454 10531 24506
rect 10583 24454 10595 24506
rect 10647 24454 10659 24506
rect 10711 24454 16705 24506
rect 16757 24454 16769 24506
rect 16821 24454 16833 24506
rect 16885 24454 16897 24506
rect 16949 24454 16961 24506
rect 17013 24454 23007 24506
rect 23059 24454 23071 24506
rect 23123 24454 23135 24506
rect 23187 24454 23199 24506
rect 23251 24454 23263 24506
rect 23315 24454 26312 24506
rect 1104 24432 26312 24454
rect 6454 24352 6460 24404
rect 6512 24392 6518 24404
rect 7561 24395 7619 24401
rect 7561 24392 7573 24395
rect 6512 24364 7573 24392
rect 6512 24352 6518 24364
rect 7561 24361 7573 24364
rect 7607 24361 7619 24395
rect 7561 24355 7619 24361
rect 8018 24352 8024 24404
rect 8076 24392 8082 24404
rect 8570 24392 8576 24404
rect 8076 24364 8576 24392
rect 8076 24352 8082 24364
rect 8570 24352 8576 24364
rect 8628 24352 8634 24404
rect 8757 24395 8815 24401
rect 8757 24361 8769 24395
rect 8803 24392 8815 24395
rect 9306 24392 9312 24404
rect 8803 24364 9312 24392
rect 8803 24361 8815 24364
rect 8757 24355 8815 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 14642 24352 14648 24404
rect 14700 24352 14706 24404
rect 14918 24352 14924 24404
rect 14976 24392 14982 24404
rect 15013 24395 15071 24401
rect 15013 24392 15025 24395
rect 14976 24364 15025 24392
rect 14976 24352 14982 24364
rect 15013 24361 15025 24364
rect 15059 24361 15071 24395
rect 15013 24355 15071 24361
rect 15105 24395 15163 24401
rect 15105 24361 15117 24395
rect 15151 24392 15163 24395
rect 15194 24392 15200 24404
rect 15151 24364 15200 24392
rect 15151 24361 15163 24364
rect 15105 24355 15163 24361
rect 15194 24352 15200 24364
rect 15252 24352 15258 24404
rect 15565 24395 15623 24401
rect 15565 24361 15577 24395
rect 15611 24361 15623 24395
rect 15565 24355 15623 24361
rect 8202 24324 8208 24336
rect 7852 24296 8208 24324
rect 5629 24259 5687 24265
rect 5629 24225 5641 24259
rect 5675 24256 5687 24259
rect 6546 24256 6552 24268
rect 5675 24228 6552 24256
rect 5675 24225 5687 24228
rect 5629 24219 5687 24225
rect 6546 24216 6552 24228
rect 6604 24216 6610 24268
rect 7762 24201 7820 24207
rect 5994 24148 6000 24200
rect 6052 24148 6058 24200
rect 7762 24167 7774 24201
rect 7808 24198 7820 24201
rect 7852 24198 7880 24296
rect 8202 24284 8208 24296
rect 8260 24284 8266 24336
rect 8846 24284 8852 24336
rect 8904 24324 8910 24336
rect 13863 24327 13921 24333
rect 8904 24296 9674 24324
rect 8904 24284 8910 24296
rect 9030 24256 9036 24268
rect 8036 24228 9036 24256
rect 8036 24198 8064 24228
rect 9030 24216 9036 24228
rect 9088 24256 9094 24268
rect 9088 24228 9536 24256
rect 9088 24216 9094 24228
rect 7808 24170 7880 24198
rect 7944 24197 8064 24198
rect 7929 24191 8064 24197
rect 7808 24167 7820 24170
rect 7762 24161 7820 24167
rect 7929 24157 7941 24191
rect 7975 24170 8064 24191
rect 7975 24157 7987 24170
rect 7929 24151 7987 24157
rect 8202 24148 8208 24200
rect 8260 24148 8266 24200
rect 8846 24188 8852 24200
rect 8312 24160 8852 24188
rect 6546 24080 6552 24132
rect 6604 24080 6610 24132
rect 7837 24123 7895 24129
rect 7837 24120 7849 24123
rect 7760 24092 7849 24120
rect 7760 24064 7788 24092
rect 7837 24089 7849 24092
rect 7883 24089 7895 24123
rect 7837 24083 7895 24089
rect 8067 24123 8125 24129
rect 8067 24089 8079 24123
rect 8113 24120 8125 24123
rect 8312 24120 8340 24160
rect 8846 24148 8852 24160
rect 8904 24148 8910 24200
rect 9125 24191 9183 24197
rect 9125 24157 9137 24191
rect 9171 24188 9183 24191
rect 9306 24188 9312 24200
rect 9171 24160 9312 24188
rect 9171 24157 9183 24160
rect 9125 24151 9183 24157
rect 9306 24148 9312 24160
rect 9364 24148 9370 24200
rect 9398 24148 9404 24200
rect 9456 24148 9462 24200
rect 9508 24197 9536 24228
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24157 9551 24191
rect 9646 24188 9674 24296
rect 13863 24293 13875 24327
rect 13909 24324 13921 24327
rect 13909 24296 14688 24324
rect 13909 24293 13921 24296
rect 13863 24287 13921 24293
rect 14660 24268 14688 24296
rect 14734 24284 14740 24336
rect 14792 24324 14798 24336
rect 15580 24324 15608 24355
rect 15746 24352 15752 24404
rect 15804 24352 15810 24404
rect 15933 24395 15991 24401
rect 15933 24361 15945 24395
rect 15979 24392 15991 24395
rect 16022 24392 16028 24404
rect 15979 24364 16028 24392
rect 15979 24361 15991 24364
rect 15933 24355 15991 24361
rect 16022 24352 16028 24364
rect 16080 24352 16086 24404
rect 16390 24352 16396 24404
rect 16448 24352 16454 24404
rect 16574 24352 16580 24404
rect 16632 24392 16638 24404
rect 17313 24395 17371 24401
rect 17313 24392 17325 24395
rect 16632 24364 17325 24392
rect 16632 24352 16638 24364
rect 17313 24361 17325 24364
rect 17359 24392 17371 24395
rect 17954 24392 17960 24404
rect 17359 24364 17960 24392
rect 17359 24361 17371 24364
rect 17313 24355 17371 24361
rect 17954 24352 17960 24364
rect 18012 24352 18018 24404
rect 20625 24395 20683 24401
rect 20625 24392 20637 24395
rect 20456 24364 20637 24392
rect 16408 24324 16436 24352
rect 17034 24324 17040 24336
rect 14792 24296 16344 24324
rect 16408 24296 17040 24324
rect 14792 24284 14798 24296
rect 10226 24216 10232 24268
rect 10284 24256 10290 24268
rect 10284 24228 11928 24256
rect 10284 24216 10290 24228
rect 11900 24200 11928 24228
rect 12434 24216 12440 24268
rect 12492 24216 12498 24268
rect 13630 24216 13636 24268
rect 13688 24256 13694 24268
rect 14185 24259 14243 24265
rect 14185 24256 14197 24259
rect 13688 24228 14197 24256
rect 13688 24216 13694 24228
rect 14185 24225 14197 24228
rect 14231 24225 14243 24259
rect 14185 24219 14243 24225
rect 14642 24216 14648 24268
rect 14700 24256 14706 24268
rect 14875 24259 14933 24265
rect 14875 24256 14887 24259
rect 14700 24228 14887 24256
rect 14700 24216 14706 24228
rect 14875 24225 14887 24228
rect 14921 24225 14933 24259
rect 14875 24219 14933 24225
rect 15473 24259 15531 24265
rect 15473 24225 15485 24259
rect 15519 24256 15531 24259
rect 15654 24256 15660 24268
rect 15519 24228 15660 24256
rect 15519 24225 15531 24228
rect 15473 24219 15531 24225
rect 15654 24216 15660 24228
rect 15712 24216 15718 24268
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24225 16267 24259
rect 16209 24219 16267 24225
rect 9769 24191 9827 24197
rect 9769 24188 9781 24191
rect 9646 24160 9781 24188
rect 9493 24151 9551 24157
rect 9769 24157 9781 24160
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 9858 24148 9864 24200
rect 9916 24148 9922 24200
rect 11606 24148 11612 24200
rect 11664 24148 11670 24200
rect 11882 24148 11888 24200
rect 11940 24188 11946 24200
rect 12069 24191 12127 24197
rect 12069 24188 12081 24191
rect 11940 24160 12081 24188
rect 11940 24148 11946 24160
rect 12069 24157 12081 24160
rect 12115 24157 12127 24191
rect 12069 24151 12127 24157
rect 13814 24148 13820 24200
rect 13872 24188 13878 24200
rect 13998 24188 14004 24200
rect 13872 24160 14004 24188
rect 13872 24148 13878 24160
rect 13998 24148 14004 24160
rect 14056 24188 14062 24200
rect 14277 24191 14335 24197
rect 14277 24188 14289 24191
rect 14056 24160 14289 24188
rect 14056 24148 14062 24160
rect 14277 24157 14289 24160
rect 14323 24188 14335 24191
rect 14734 24188 14740 24200
rect 14323 24160 14740 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 14734 24148 14740 24160
rect 14792 24148 14798 24200
rect 15197 24191 15255 24197
rect 15197 24157 15209 24191
rect 15243 24188 15255 24191
rect 15243 24160 15424 24188
rect 15243 24157 15255 24160
rect 15197 24151 15255 24157
rect 8113 24092 8340 24120
rect 8113 24089 8125 24092
rect 8067 24083 8125 24089
rect 8386 24080 8392 24132
rect 8444 24080 8450 24132
rect 8478 24080 8484 24132
rect 8536 24120 8542 24132
rect 8941 24123 8999 24129
rect 8536 24092 8892 24120
rect 8536 24080 8542 24092
rect 7423 24055 7481 24061
rect 7423 24021 7435 24055
rect 7469 24052 7481 24055
rect 7650 24052 7656 24064
rect 7469 24024 7656 24052
rect 7469 24021 7481 24024
rect 7423 24015 7481 24021
rect 7650 24012 7656 24024
rect 7708 24012 7714 24064
rect 7742 24012 7748 24064
rect 7800 24012 7806 24064
rect 8294 24012 8300 24064
rect 8352 24052 8358 24064
rect 8589 24055 8647 24061
rect 8589 24052 8601 24055
rect 8352 24024 8601 24052
rect 8352 24012 8358 24024
rect 8589 24021 8601 24024
rect 8635 24021 8647 24055
rect 8864 24052 8892 24092
rect 8941 24089 8953 24123
rect 8987 24120 8999 24123
rect 9677 24123 9735 24129
rect 9677 24120 9689 24123
rect 8987 24092 9689 24120
rect 8987 24089 8999 24092
rect 8941 24083 8999 24089
rect 9677 24089 9689 24092
rect 9723 24089 9735 24123
rect 9677 24083 9735 24089
rect 10505 24123 10563 24129
rect 10505 24089 10517 24123
rect 10551 24089 10563 24123
rect 10505 24083 10563 24089
rect 9309 24055 9367 24061
rect 9309 24052 9321 24055
rect 8864 24024 9321 24052
rect 8589 24015 8647 24021
rect 9309 24021 9321 24024
rect 9355 24021 9367 24055
rect 9309 24015 9367 24021
rect 9490 24012 9496 24064
rect 9548 24052 9554 24064
rect 9950 24052 9956 24064
rect 9548 24024 9956 24052
rect 9548 24012 9554 24024
rect 9950 24012 9956 24024
rect 10008 24012 10014 24064
rect 10045 24055 10103 24061
rect 10045 24021 10057 24055
rect 10091 24052 10103 24055
rect 10520 24052 10548 24083
rect 12986 24080 12992 24132
rect 13044 24080 13050 24132
rect 15286 24080 15292 24132
rect 15344 24080 15350 24132
rect 15396 24120 15424 24160
rect 15562 24148 15568 24200
rect 15620 24148 15626 24200
rect 16117 24191 16175 24197
rect 16117 24188 16129 24191
rect 15672 24160 16129 24188
rect 15580 24120 15608 24148
rect 15396 24092 15608 24120
rect 10091 24024 10548 24052
rect 11977 24055 12035 24061
rect 10091 24021 10103 24024
rect 10045 24015 10103 24021
rect 11977 24021 11989 24055
rect 12023 24052 12035 24055
rect 12066 24052 12072 24064
rect 12023 24024 12072 24052
rect 12023 24021 12035 24024
rect 11977 24015 12035 24021
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 15304 24052 15332 24080
rect 15672 24052 15700 24160
rect 16117 24157 16129 24160
rect 16163 24157 16175 24191
rect 16117 24151 16175 24157
rect 15746 24080 15752 24132
rect 15804 24120 15810 24132
rect 16224 24120 16252 24219
rect 16316 24197 16344 24296
rect 17034 24284 17040 24296
rect 17092 24284 17098 24336
rect 17218 24284 17224 24336
rect 17276 24324 17282 24336
rect 17773 24327 17831 24333
rect 17773 24324 17785 24327
rect 17276 24296 17785 24324
rect 17276 24284 17282 24296
rect 17773 24293 17785 24296
rect 17819 24293 17831 24327
rect 17773 24287 17831 24293
rect 16390 24216 16396 24268
rect 16448 24216 16454 24268
rect 17494 24216 17500 24268
rect 17552 24216 17558 24268
rect 20456 24256 20484 24364
rect 20625 24361 20637 24364
rect 20671 24361 20683 24395
rect 20625 24355 20683 24361
rect 20714 24352 20720 24404
rect 20772 24392 20778 24404
rect 21085 24395 21143 24401
rect 21085 24392 21097 24395
rect 20772 24364 21097 24392
rect 20772 24352 20778 24364
rect 21085 24361 21097 24364
rect 21131 24361 21143 24395
rect 21085 24355 21143 24361
rect 21174 24352 21180 24404
rect 21232 24392 21238 24404
rect 22370 24392 22376 24404
rect 21232 24364 22376 24392
rect 21232 24352 21238 24364
rect 22370 24352 22376 24364
rect 22428 24352 22434 24404
rect 22465 24395 22523 24401
rect 22465 24361 22477 24395
rect 22511 24392 22523 24395
rect 22554 24392 22560 24404
rect 22511 24364 22560 24392
rect 22511 24361 22523 24364
rect 22465 24355 22523 24361
rect 22554 24352 22560 24364
rect 22612 24352 22618 24404
rect 23382 24352 23388 24404
rect 23440 24392 23446 24404
rect 23440 24364 24072 24392
rect 23440 24352 23446 24364
rect 20530 24284 20536 24336
rect 20588 24324 20594 24336
rect 23474 24324 23480 24336
rect 20588 24296 23480 24324
rect 20588 24284 20594 24296
rect 23474 24284 23480 24296
rect 23532 24284 23538 24336
rect 23753 24327 23811 24333
rect 23753 24293 23765 24327
rect 23799 24293 23811 24327
rect 23753 24287 23811 24293
rect 20809 24259 20867 24265
rect 20456 24228 20760 24256
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24188 16359 24191
rect 16482 24188 16488 24200
rect 16347 24160 16488 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 17034 24148 17040 24200
rect 17092 24188 17098 24200
rect 17221 24191 17279 24197
rect 17221 24188 17233 24191
rect 17092 24160 17233 24188
rect 17092 24148 17098 24160
rect 17221 24157 17233 24160
rect 17267 24188 17279 24191
rect 18138 24188 18144 24200
rect 17267 24160 18144 24188
rect 17267 24157 17279 24160
rect 17221 24151 17279 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18874 24148 18880 24200
rect 18932 24188 18938 24200
rect 20070 24188 20076 24200
rect 18932 24160 20076 24188
rect 18932 24148 18938 24160
rect 20070 24148 20076 24160
rect 20128 24188 20134 24200
rect 20533 24191 20591 24197
rect 20533 24188 20545 24191
rect 20128 24160 20545 24188
rect 20128 24148 20134 24160
rect 20533 24157 20545 24160
rect 20579 24157 20591 24191
rect 20732 24188 20760 24228
rect 20809 24225 20821 24259
rect 20855 24256 20867 24259
rect 20898 24256 20904 24268
rect 20855 24228 20904 24256
rect 20855 24225 20867 24228
rect 20809 24219 20867 24225
rect 20898 24216 20904 24228
rect 20956 24256 20962 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 20956 24228 21281 24256
rect 20956 24216 20962 24228
rect 21269 24225 21281 24228
rect 21315 24225 21327 24259
rect 21269 24219 21327 24225
rect 22186 24216 22192 24268
rect 22244 24256 22250 24268
rect 23768 24256 23796 24287
rect 22244 24228 23796 24256
rect 22244 24216 22250 24228
rect 21082 24188 21088 24200
rect 20732 24160 21088 24188
rect 20533 24151 20591 24157
rect 15804 24092 16252 24120
rect 20548 24120 20576 24151
rect 21082 24148 21088 24160
rect 21140 24148 21146 24200
rect 21177 24191 21235 24197
rect 21177 24157 21189 24191
rect 21223 24188 21235 24191
rect 21358 24188 21364 24200
rect 21223 24160 21364 24188
rect 21223 24157 21235 24160
rect 21177 24151 21235 24157
rect 21358 24148 21364 24160
rect 21416 24148 21422 24200
rect 22278 24148 22284 24200
rect 22336 24188 22342 24200
rect 22465 24191 22523 24197
rect 22465 24188 22477 24191
rect 22336 24160 22477 24188
rect 22336 24148 22342 24160
rect 22465 24157 22477 24160
rect 22511 24157 22523 24191
rect 22465 24151 22523 24157
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 20714 24120 20720 24132
rect 20548 24092 20720 24120
rect 15804 24080 15810 24092
rect 20714 24080 20720 24092
rect 20772 24080 20778 24132
rect 20806 24080 20812 24132
rect 20864 24120 20870 24132
rect 22664 24120 22692 24151
rect 23106 24148 23112 24200
rect 23164 24148 23170 24200
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 23566 24188 23572 24200
rect 23523 24160 23572 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 24044 24197 24072 24364
rect 23937 24191 23995 24197
rect 23937 24188 23949 24191
rect 23676 24160 23949 24188
rect 20864 24092 22692 24120
rect 20864 24080 20870 24092
rect 15304 24024 15700 24052
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 21358 24052 21364 24064
rect 19944 24024 21364 24052
rect 19944 24012 19950 24024
rect 21358 24012 21364 24024
rect 21416 24012 21422 24064
rect 22664 24052 22692 24092
rect 22922 24080 22928 24132
rect 22980 24120 22986 24132
rect 23293 24123 23351 24129
rect 23293 24120 23305 24123
rect 22980 24092 23305 24120
rect 22980 24080 22986 24092
rect 23293 24089 23305 24092
rect 23339 24089 23351 24123
rect 23293 24083 23351 24089
rect 23385 24123 23443 24129
rect 23385 24089 23397 24123
rect 23431 24120 23443 24123
rect 23676 24120 23704 24160
rect 23937 24157 23949 24160
rect 23983 24157 23995 24191
rect 23937 24151 23995 24157
rect 24029 24191 24087 24197
rect 24029 24157 24041 24191
rect 24075 24157 24087 24191
rect 24029 24151 24087 24157
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 24360 24160 24409 24188
rect 24360 24148 24366 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24397 24151 24455 24157
rect 23431 24092 23704 24120
rect 23431 24089 23443 24092
rect 23385 24083 23443 24089
rect 23400 24052 23428 24083
rect 23750 24080 23756 24132
rect 23808 24120 23814 24132
rect 25038 24120 25044 24132
rect 23808 24092 25044 24120
rect 23808 24080 23814 24092
rect 25038 24080 25044 24092
rect 25096 24080 25102 24132
rect 22664 24024 23428 24052
rect 23474 24012 23480 24064
rect 23532 24052 23538 24064
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23532 24024 23673 24052
rect 23532 24012 23538 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 24486 24012 24492 24064
rect 24544 24012 24550 24064
rect 1104 23962 26312 23984
rect 1104 23910 4761 23962
rect 4813 23910 4825 23962
rect 4877 23910 4889 23962
rect 4941 23910 4953 23962
rect 5005 23910 5017 23962
rect 5069 23910 11063 23962
rect 11115 23910 11127 23962
rect 11179 23910 11191 23962
rect 11243 23910 11255 23962
rect 11307 23910 11319 23962
rect 11371 23910 17365 23962
rect 17417 23910 17429 23962
rect 17481 23910 17493 23962
rect 17545 23910 17557 23962
rect 17609 23910 17621 23962
rect 17673 23910 23667 23962
rect 23719 23910 23731 23962
rect 23783 23910 23795 23962
rect 23847 23910 23859 23962
rect 23911 23910 23923 23962
rect 23975 23910 26312 23962
rect 1104 23888 26312 23910
rect 6546 23808 6552 23860
rect 6604 23808 6610 23860
rect 6825 23851 6883 23857
rect 6825 23817 6837 23851
rect 6871 23817 6883 23851
rect 6825 23811 6883 23817
rect 3694 23740 3700 23792
rect 3752 23780 3758 23792
rect 4249 23783 4307 23789
rect 4249 23780 4261 23783
rect 3752 23752 4261 23780
rect 3752 23740 3758 23752
rect 4249 23749 4261 23752
rect 4295 23749 4307 23783
rect 4249 23743 4307 23749
rect 4433 23783 4491 23789
rect 4433 23749 4445 23783
rect 4479 23780 4491 23783
rect 5166 23780 5172 23792
rect 4479 23752 5172 23780
rect 4479 23749 4491 23752
rect 4433 23743 4491 23749
rect 5166 23740 5172 23752
rect 5224 23740 5230 23792
rect 5994 23740 6000 23792
rect 6052 23780 6058 23792
rect 6840 23780 6868 23811
rect 7742 23808 7748 23860
rect 7800 23848 7806 23860
rect 8297 23851 8355 23857
rect 8297 23848 8309 23851
rect 7800 23820 8309 23848
rect 7800 23808 7806 23820
rect 8297 23817 8309 23820
rect 8343 23817 8355 23851
rect 8297 23811 8355 23817
rect 8481 23851 8539 23857
rect 8481 23817 8493 23851
rect 8527 23848 8539 23851
rect 8846 23848 8852 23860
rect 8527 23820 8852 23848
rect 8527 23817 8539 23820
rect 8481 23811 8539 23817
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9398 23808 9404 23860
rect 9456 23848 9462 23860
rect 10413 23851 10471 23857
rect 10413 23848 10425 23851
rect 9456 23820 10425 23848
rect 9456 23808 9462 23820
rect 10413 23817 10425 23820
rect 10459 23817 10471 23851
rect 10413 23811 10471 23817
rect 11606 23808 11612 23860
rect 11664 23808 11670 23860
rect 12986 23808 12992 23860
rect 13044 23848 13050 23860
rect 13081 23851 13139 23857
rect 13081 23848 13093 23851
rect 13044 23820 13093 23848
rect 13044 23808 13050 23820
rect 13081 23817 13093 23820
rect 13127 23817 13139 23851
rect 13081 23811 13139 23817
rect 13630 23808 13636 23860
rect 13688 23848 13694 23860
rect 15013 23851 15071 23857
rect 15013 23848 15025 23851
rect 13688 23820 15025 23848
rect 13688 23808 13694 23820
rect 15013 23817 15025 23820
rect 15059 23848 15071 23851
rect 15765 23851 15823 23857
rect 15765 23848 15777 23851
rect 15059 23820 15777 23848
rect 15059 23817 15071 23820
rect 15013 23811 15071 23817
rect 15765 23817 15777 23820
rect 15811 23817 15823 23851
rect 15765 23811 15823 23817
rect 15933 23851 15991 23857
rect 15933 23817 15945 23851
rect 15979 23848 15991 23851
rect 16574 23848 16580 23860
rect 15979 23820 16580 23848
rect 15979 23817 15991 23820
rect 15933 23811 15991 23817
rect 16574 23808 16580 23820
rect 16632 23808 16638 23860
rect 20898 23808 20904 23860
rect 20956 23808 20962 23860
rect 22373 23851 22431 23857
rect 22373 23817 22385 23851
rect 22419 23848 22431 23851
rect 22554 23848 22560 23860
rect 22419 23820 22560 23848
rect 22419 23817 22431 23820
rect 22373 23811 22431 23817
rect 22554 23808 22560 23820
rect 22612 23808 22618 23860
rect 22922 23808 22928 23860
rect 22980 23808 22986 23860
rect 7834 23780 7840 23792
rect 6052 23752 6868 23780
rect 7024 23752 7840 23780
rect 6052 23740 6058 23752
rect 5353 23715 5411 23721
rect 5353 23712 5365 23715
rect 4724 23684 5365 23712
rect 4157 23647 4215 23653
rect 4157 23613 4169 23647
rect 4203 23613 4215 23647
rect 4157 23607 4215 23613
rect 3694 23468 3700 23520
rect 3752 23468 3758 23520
rect 4172 23508 4200 23607
rect 4724 23585 4752 23684
rect 5353 23681 5365 23684
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 6454 23672 6460 23724
rect 6512 23672 6518 23724
rect 7024 23721 7052 23752
rect 7834 23740 7840 23752
rect 7892 23740 7898 23792
rect 8202 23780 8208 23792
rect 8036 23752 8208 23780
rect 7009 23715 7067 23721
rect 7009 23681 7021 23715
rect 7055 23681 7067 23715
rect 7009 23675 7067 23681
rect 7282 23672 7288 23724
rect 7340 23672 7346 23724
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 7484 23684 7757 23712
rect 7101 23647 7159 23653
rect 7101 23613 7113 23647
rect 7147 23613 7159 23647
rect 7101 23607 7159 23613
rect 7193 23647 7251 23653
rect 7193 23613 7205 23647
rect 7239 23644 7251 23647
rect 7484 23644 7512 23684
rect 7745 23681 7757 23684
rect 7791 23712 7803 23715
rect 8036 23712 8064 23752
rect 8202 23740 8208 23752
rect 8260 23740 8266 23792
rect 9306 23780 9312 23792
rect 8588 23752 9312 23780
rect 7791 23684 8064 23712
rect 8113 23715 8171 23721
rect 7791 23681 7803 23684
rect 7745 23675 7803 23681
rect 8113 23681 8125 23715
rect 8159 23712 8171 23715
rect 8478 23712 8484 23724
rect 8159 23684 8484 23712
rect 8159 23681 8171 23684
rect 8113 23675 8171 23681
rect 8478 23672 8484 23684
rect 8536 23672 8542 23724
rect 7239 23616 7512 23644
rect 7239 23613 7251 23616
rect 7193 23607 7251 23613
rect 4709 23579 4767 23585
rect 4709 23545 4721 23579
rect 4755 23545 4767 23579
rect 4709 23539 4767 23545
rect 5534 23536 5540 23588
rect 5592 23536 5598 23588
rect 7116 23576 7144 23607
rect 7558 23604 7564 23656
rect 7616 23644 7622 23656
rect 8588 23644 8616 23752
rect 8864 23721 8892 23752
rect 9306 23740 9312 23752
rect 9364 23740 9370 23792
rect 9582 23740 9588 23792
rect 9640 23740 9646 23792
rect 9794 23783 9852 23789
rect 9794 23749 9806 23783
rect 9840 23780 9852 23783
rect 10134 23780 10140 23792
rect 9840 23752 10140 23780
rect 9840 23749 9852 23752
rect 9794 23743 9852 23749
rect 10134 23740 10140 23752
rect 10192 23740 10198 23792
rect 14918 23780 14924 23792
rect 14292 23752 14924 23780
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23681 8723 23715
rect 8665 23675 8723 23681
rect 8849 23715 8907 23721
rect 8849 23681 8861 23715
rect 8895 23681 8907 23715
rect 8849 23675 8907 23681
rect 7616 23616 8616 23644
rect 8680 23644 8708 23675
rect 8938 23672 8944 23724
rect 8996 23672 9002 23724
rect 9214 23672 9220 23724
rect 9272 23672 9278 23724
rect 9490 23672 9496 23724
rect 9548 23672 9554 23724
rect 9600 23712 9628 23740
rect 9677 23721 9735 23727
rect 14292 23724 14320 23752
rect 9677 23712 9689 23721
rect 9600 23687 9689 23712
rect 9723 23687 9735 23721
rect 9600 23684 9735 23687
rect 9677 23681 9735 23684
rect 9950 23672 9956 23724
rect 10008 23672 10014 23724
rect 10045 23715 10103 23721
rect 10045 23681 10057 23715
rect 10091 23712 10103 23715
rect 10318 23712 10324 23724
rect 10091 23684 10324 23712
rect 10091 23681 10103 23684
rect 10045 23675 10103 23681
rect 10318 23672 10324 23684
rect 10376 23712 10382 23724
rect 10376 23684 10916 23712
rect 10376 23672 10382 23684
rect 9030 23644 9036 23656
rect 8680 23616 9036 23644
rect 7616 23604 7622 23616
rect 7466 23576 7472 23588
rect 7116 23548 7472 23576
rect 7466 23536 7472 23548
rect 7524 23536 7530 23588
rect 7650 23536 7656 23588
rect 7708 23576 7714 23588
rect 8386 23576 8392 23588
rect 7708 23548 8392 23576
rect 7708 23536 7714 23548
rect 5626 23508 5632 23520
rect 4172 23480 5632 23508
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 8128 23517 8156 23548
rect 8386 23536 8392 23548
rect 8444 23576 8450 23588
rect 8680 23576 8708 23616
rect 9030 23604 9036 23616
rect 9088 23604 9094 23656
rect 8444 23548 8708 23576
rect 8444 23536 8450 23548
rect 8754 23536 8760 23588
rect 8812 23585 8818 23588
rect 8812 23576 8819 23585
rect 9122 23576 9128 23588
rect 8812 23548 9128 23576
rect 8812 23539 8819 23548
rect 8812 23536 8818 23539
rect 9122 23536 9128 23548
rect 9180 23536 9186 23588
rect 8113 23511 8171 23517
rect 8113 23477 8125 23511
rect 8159 23477 8171 23511
rect 8113 23471 8171 23477
rect 8202 23468 8208 23520
rect 8260 23508 8266 23520
rect 8772 23508 8800 23536
rect 8260 23480 8800 23508
rect 9232 23508 9260 23672
rect 9355 23647 9413 23653
rect 9355 23613 9367 23647
rect 9401 23644 9413 23647
rect 9508 23644 9536 23672
rect 9401 23616 9536 23644
rect 9401 23613 9413 23616
rect 9355 23607 9413 23613
rect 9582 23604 9588 23656
rect 9640 23604 9646 23656
rect 10597 23647 10655 23653
rect 10597 23613 10609 23647
rect 10643 23613 10655 23647
rect 10597 23607 10655 23613
rect 9490 23536 9496 23588
rect 9548 23536 9554 23588
rect 10134 23536 10140 23588
rect 10192 23576 10198 23588
rect 10612 23576 10640 23607
rect 10686 23604 10692 23656
rect 10744 23604 10750 23656
rect 10778 23604 10784 23656
rect 10836 23604 10842 23656
rect 10888 23653 10916 23684
rect 11054 23672 11060 23724
rect 11112 23712 11118 23724
rect 11517 23715 11575 23721
rect 11517 23712 11529 23715
rect 11112 23684 11529 23712
rect 11112 23672 11118 23684
rect 11517 23681 11529 23684
rect 11563 23712 11575 23715
rect 12894 23712 12900 23724
rect 11563 23684 12900 23712
rect 11563 23681 11575 23684
rect 11517 23675 11575 23681
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 12989 23715 13047 23721
rect 12989 23681 13001 23715
rect 13035 23712 13047 23715
rect 13722 23712 13728 23724
rect 13035 23684 13728 23712
rect 13035 23681 13047 23684
rect 12989 23675 13047 23681
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 13814 23672 13820 23724
rect 13872 23672 13878 23724
rect 14274 23672 14280 23724
rect 14332 23672 14338 23724
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23712 14519 23715
rect 14642 23712 14648 23724
rect 14507 23684 14648 23712
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 14642 23672 14648 23684
rect 14700 23712 14706 23724
rect 14844 23721 14872 23752
rect 14918 23740 14924 23752
rect 14976 23780 14982 23792
rect 15286 23780 15292 23792
rect 14976 23752 15292 23780
rect 14976 23740 14982 23752
rect 15286 23740 15292 23752
rect 15344 23740 15350 23792
rect 15562 23740 15568 23792
rect 15620 23780 15626 23792
rect 16298 23780 16304 23792
rect 15620 23752 16304 23780
rect 15620 23740 15626 23752
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 21085 23783 21143 23789
rect 21085 23749 21097 23783
rect 21131 23780 21143 23783
rect 21174 23780 21180 23792
rect 21131 23752 21180 23780
rect 21131 23749 21143 23752
rect 21085 23743 21143 23749
rect 21174 23740 21180 23752
rect 21232 23740 21238 23792
rect 21358 23789 21364 23792
rect 21301 23783 21364 23789
rect 21301 23749 21313 23783
rect 21347 23749 21364 23783
rect 21301 23743 21364 23749
rect 21358 23740 21364 23743
rect 21416 23740 21422 23792
rect 22278 23780 22284 23792
rect 22066 23752 22284 23780
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 14700 23684 14749 23712
rect 14700 23672 14706 23684
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 20717 23715 20775 23721
rect 20717 23681 20729 23715
rect 20763 23681 20775 23715
rect 20717 23675 20775 23681
rect 10873 23647 10931 23653
rect 10873 23613 10885 23647
rect 10919 23644 10931 23647
rect 12066 23644 12072 23656
rect 10919 23616 12072 23644
rect 10919 23613 10931 23616
rect 10873 23607 10931 23613
rect 12066 23604 12072 23616
rect 12124 23604 12130 23656
rect 13906 23604 13912 23656
rect 13964 23644 13970 23656
rect 14369 23647 14427 23653
rect 14369 23644 14381 23647
rect 13964 23616 14381 23644
rect 13964 23604 13970 23616
rect 14369 23613 14381 23616
rect 14415 23613 14427 23647
rect 14752 23644 14780 23675
rect 15654 23644 15660 23656
rect 14752 23616 15660 23644
rect 14369 23607 14427 23613
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 20732 23644 20760 23675
rect 20990 23672 20996 23724
rect 21048 23672 21054 23724
rect 20732 23616 21496 23644
rect 12802 23576 12808 23588
rect 10192 23548 12808 23576
rect 10192 23536 10198 23548
rect 12802 23536 12808 23548
rect 12860 23536 12866 23588
rect 14185 23579 14243 23585
rect 14185 23545 14197 23579
rect 14231 23576 14243 23579
rect 14458 23576 14464 23588
rect 14231 23548 14464 23576
rect 14231 23545 14243 23548
rect 14185 23539 14243 23545
rect 14458 23536 14464 23548
rect 14516 23536 14522 23588
rect 21468 23585 21496 23616
rect 21453 23579 21511 23585
rect 21453 23545 21465 23579
rect 21499 23576 21511 23579
rect 22066 23576 22094 23752
rect 22278 23740 22284 23752
rect 22336 23780 22342 23792
rect 22741 23783 22799 23789
rect 22741 23780 22753 23783
rect 22336 23752 22753 23780
rect 22336 23740 22342 23752
rect 22741 23749 22753 23752
rect 22787 23749 22799 23783
rect 24486 23780 24492 23792
rect 24426 23752 24492 23780
rect 22741 23743 22799 23749
rect 24486 23740 24492 23752
rect 24544 23740 24550 23792
rect 22186 23672 22192 23724
rect 22244 23672 22250 23724
rect 22465 23715 22523 23721
rect 22465 23681 22477 23715
rect 22511 23681 22523 23715
rect 22465 23675 22523 23681
rect 21499 23548 22094 23576
rect 22480 23576 22508 23675
rect 22554 23672 22560 23724
rect 22612 23672 22618 23724
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23712 23443 23715
rect 23474 23712 23480 23724
rect 23431 23684 23480 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 22646 23604 22652 23656
rect 22704 23644 22710 23656
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22704 23616 23029 23644
rect 22704 23604 22710 23616
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 23017 23607 23075 23613
rect 22480 23548 23060 23576
rect 21499 23545 21511 23548
rect 21453 23539 21511 23545
rect 9950 23508 9956 23520
rect 9232 23480 9956 23508
rect 8260 23468 8266 23480
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 10042 23468 10048 23520
rect 10100 23508 10106 23520
rect 10229 23511 10287 23517
rect 10229 23508 10241 23511
rect 10100 23480 10241 23508
rect 10100 23468 10106 23480
rect 10229 23477 10241 23480
rect 10275 23477 10287 23511
rect 10229 23471 10287 23477
rect 10686 23468 10692 23520
rect 10744 23508 10750 23520
rect 11698 23508 11704 23520
rect 10744 23480 11704 23508
rect 10744 23468 10750 23480
rect 11698 23468 11704 23480
rect 11756 23468 11762 23520
rect 15749 23511 15807 23517
rect 15749 23477 15761 23511
rect 15795 23508 15807 23511
rect 16482 23508 16488 23520
rect 15795 23480 16488 23508
rect 15795 23477 15807 23480
rect 15749 23471 15807 23477
rect 16482 23468 16488 23480
rect 16540 23508 16546 23520
rect 17034 23508 17040 23520
rect 16540 23480 17040 23508
rect 16540 23468 16546 23480
rect 17034 23468 17040 23480
rect 17092 23468 17098 23520
rect 20438 23468 20444 23520
rect 20496 23508 20502 23520
rect 20533 23511 20591 23517
rect 20533 23508 20545 23511
rect 20496 23480 20545 23508
rect 20496 23468 20502 23480
rect 20533 23477 20545 23480
rect 20579 23477 20591 23511
rect 20533 23471 20591 23477
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 21266 23508 21272 23520
rect 20772 23480 21272 23508
rect 20772 23468 20778 23480
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 22922 23508 22928 23520
rect 22235 23480 22928 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 23032 23508 23060 23548
rect 23382 23508 23388 23520
rect 23032 23480 23388 23508
rect 23382 23468 23388 23480
rect 23440 23468 23446 23520
rect 23658 23468 23664 23520
rect 23716 23508 23722 23520
rect 24765 23511 24823 23517
rect 24765 23508 24777 23511
rect 23716 23480 24777 23508
rect 23716 23468 23722 23480
rect 24765 23477 24777 23480
rect 24811 23477 24823 23511
rect 24765 23471 24823 23477
rect 1104 23418 26312 23440
rect 1104 23366 4101 23418
rect 4153 23366 4165 23418
rect 4217 23366 4229 23418
rect 4281 23366 4293 23418
rect 4345 23366 4357 23418
rect 4409 23366 10403 23418
rect 10455 23366 10467 23418
rect 10519 23366 10531 23418
rect 10583 23366 10595 23418
rect 10647 23366 10659 23418
rect 10711 23366 16705 23418
rect 16757 23366 16769 23418
rect 16821 23366 16833 23418
rect 16885 23366 16897 23418
rect 16949 23366 16961 23418
rect 17013 23366 23007 23418
rect 23059 23366 23071 23418
rect 23123 23366 23135 23418
rect 23187 23366 23199 23418
rect 23251 23366 23263 23418
rect 23315 23366 26312 23418
rect 1104 23344 26312 23366
rect 5537 23307 5595 23313
rect 5537 23273 5549 23307
rect 5583 23304 5595 23307
rect 5626 23304 5632 23316
rect 5583 23276 5632 23304
rect 5583 23273 5595 23276
rect 5537 23267 5595 23273
rect 5626 23264 5632 23276
rect 5684 23264 5690 23316
rect 9030 23264 9036 23316
rect 9088 23304 9094 23316
rect 9766 23304 9772 23316
rect 9088 23276 9772 23304
rect 9088 23264 9094 23276
rect 9766 23264 9772 23276
rect 9824 23264 9830 23316
rect 9858 23264 9864 23316
rect 9916 23264 9922 23316
rect 17129 23307 17187 23313
rect 17129 23273 17141 23307
rect 17175 23304 17187 23307
rect 19610 23304 19616 23316
rect 17175 23276 19616 23304
rect 17175 23273 17187 23276
rect 17129 23267 17187 23273
rect 19610 23264 19616 23276
rect 19668 23304 19674 23316
rect 20622 23304 20628 23316
rect 19668 23276 20628 23304
rect 19668 23264 19674 23276
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 20809 23307 20867 23313
rect 20809 23304 20821 23307
rect 20772 23276 20821 23304
rect 20772 23264 20778 23276
rect 20809 23273 20821 23276
rect 20855 23273 20867 23307
rect 20809 23267 20867 23273
rect 20901 23307 20959 23313
rect 20901 23273 20913 23307
rect 20947 23304 20959 23307
rect 20990 23304 20996 23316
rect 20947 23276 20996 23304
rect 20947 23273 20959 23276
rect 20901 23267 20959 23273
rect 20990 23264 20996 23276
rect 21048 23264 21054 23316
rect 21729 23307 21787 23313
rect 21729 23304 21741 23307
rect 21284 23276 21741 23304
rect 5644 23177 5672 23264
rect 9950 23196 9956 23248
rect 10008 23236 10014 23248
rect 18046 23236 18052 23248
rect 10008 23208 18052 23236
rect 10008 23196 10014 23208
rect 18046 23196 18052 23208
rect 18104 23196 18110 23248
rect 19794 23196 19800 23248
rect 19852 23236 19858 23248
rect 19852 23208 21220 23236
rect 19852 23196 19858 23208
rect 5629 23171 5687 23177
rect 5629 23137 5641 23171
rect 5675 23137 5687 23171
rect 5629 23131 5687 23137
rect 9122 23128 9128 23180
rect 9180 23168 9186 23180
rect 12986 23168 12992 23180
rect 9180 23140 12992 23168
rect 9180 23128 9186 23140
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18012 23140 18368 23168
rect 18012 23128 18018 23140
rect 3602 23060 3608 23112
rect 3660 23100 3666 23112
rect 3789 23103 3847 23109
rect 3789 23100 3801 23103
rect 3660 23072 3801 23100
rect 3660 23060 3666 23072
rect 3789 23069 3801 23072
rect 3835 23069 3847 23103
rect 3789 23063 3847 23069
rect 5994 23060 6000 23112
rect 6052 23100 6058 23112
rect 6365 23103 6423 23109
rect 6365 23100 6377 23103
rect 6052 23072 6377 23100
rect 6052 23060 6058 23072
rect 6365 23069 6377 23072
rect 6411 23069 6423 23103
rect 6365 23063 6423 23069
rect 9582 23060 9588 23112
rect 9640 23100 9646 23112
rect 9769 23103 9827 23109
rect 9769 23100 9781 23103
rect 9640 23072 9781 23100
rect 9640 23060 9646 23072
rect 9769 23069 9781 23072
rect 9815 23069 9827 23103
rect 9769 23063 9827 23069
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23100 10011 23103
rect 10042 23100 10048 23112
rect 9999 23072 10048 23100
rect 9999 23069 10011 23072
rect 9953 23063 10011 23069
rect 10042 23060 10048 23072
rect 10100 23060 10106 23112
rect 16390 23060 16396 23112
rect 16448 23100 16454 23112
rect 18340 23109 18368 23140
rect 20070 23128 20076 23180
rect 20128 23128 20134 23180
rect 20714 23168 20720 23180
rect 20640 23140 20720 23168
rect 16761 23103 16819 23109
rect 16761 23100 16773 23103
rect 16448 23072 16773 23100
rect 16448 23060 16454 23072
rect 16761 23069 16773 23072
rect 16807 23069 16819 23103
rect 16761 23063 16819 23069
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23069 18199 23103
rect 18141 23063 18199 23069
rect 18325 23103 18383 23109
rect 18325 23069 18337 23103
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23100 18475 23103
rect 18506 23100 18512 23112
rect 18463 23072 18512 23100
rect 18463 23069 18475 23072
rect 18417 23063 18475 23069
rect 4062 22992 4068 23044
rect 4120 22992 4126 23044
rect 6457 23035 6515 23041
rect 6457 23032 6469 23035
rect 5290 23004 6469 23032
rect 6457 23001 6469 23004
rect 6503 23001 6515 23035
rect 6457 22995 6515 23001
rect 15930 22992 15936 23044
rect 15988 23032 15994 23044
rect 15988 23004 17356 23032
rect 15988 22992 15994 23004
rect 6270 22924 6276 22976
rect 6328 22924 6334 22976
rect 11974 22924 11980 22976
rect 12032 22964 12038 22976
rect 16206 22964 16212 22976
rect 12032 22936 16212 22964
rect 12032 22924 12038 22936
rect 16206 22924 16212 22936
rect 16264 22924 16270 22976
rect 17126 22924 17132 22976
rect 17184 22924 17190 22976
rect 17328 22973 17356 23004
rect 17862 22992 17868 23044
rect 17920 23032 17926 23044
rect 18156 23032 18184 23063
rect 18506 23060 18512 23072
rect 18564 23060 18570 23112
rect 19702 23060 19708 23112
rect 19760 23100 19766 23112
rect 19981 23103 20039 23109
rect 19981 23100 19993 23103
rect 19760 23072 19993 23100
rect 19760 23060 19766 23072
rect 19981 23069 19993 23072
rect 20027 23069 20039 23103
rect 19981 23063 20039 23069
rect 20162 23060 20168 23112
rect 20220 23060 20226 23112
rect 20254 23062 20260 23114
rect 20312 23109 20318 23114
rect 20312 23103 20361 23109
rect 20312 23069 20315 23103
rect 20349 23102 20361 23103
rect 20349 23072 20392 23102
rect 20349 23069 20361 23072
rect 20312 23063 20361 23069
rect 20312 23062 20318 23063
rect 20438 23060 20444 23112
rect 20496 23060 20502 23112
rect 20640 23109 20668 23140
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 20990 23128 20996 23180
rect 21048 23168 21054 23180
rect 21192 23177 21220 23208
rect 21284 23180 21312 23276
rect 21729 23273 21741 23276
rect 21775 23304 21787 23307
rect 21775 23276 22324 23304
rect 21775 23273 21787 23276
rect 21729 23267 21787 23273
rect 21358 23196 21364 23248
rect 21416 23236 21422 23248
rect 21913 23239 21971 23245
rect 21913 23236 21925 23239
rect 21416 23208 21925 23236
rect 21416 23196 21422 23208
rect 21913 23205 21925 23208
rect 21959 23205 21971 23239
rect 21913 23199 21971 23205
rect 21177 23171 21235 23177
rect 21177 23168 21189 23171
rect 21048 23140 21189 23168
rect 21048 23128 21054 23140
rect 21177 23137 21189 23140
rect 21223 23137 21235 23171
rect 21177 23131 21235 23137
rect 21266 23128 21272 23180
rect 21324 23128 21330 23180
rect 22189 23171 22247 23177
rect 22189 23168 22201 23171
rect 22066 23140 22201 23168
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 20806 23060 20812 23112
rect 20864 23060 20870 23112
rect 21082 23060 21088 23112
rect 21140 23060 21146 23112
rect 21361 23103 21419 23109
rect 21361 23069 21373 23103
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 17920 23004 18368 23032
rect 17920 22992 17926 23004
rect 18340 22976 18368 23004
rect 19242 22992 19248 23044
rect 19300 23032 19306 23044
rect 19886 23032 19892 23044
rect 19300 23004 19892 23032
rect 19300 22992 19306 23004
rect 19886 22992 19892 23004
rect 19944 22992 19950 23044
rect 20533 23035 20591 23041
rect 20533 23001 20545 23035
rect 20579 23032 20591 23035
rect 20824 23032 20852 23060
rect 20579 23004 20852 23032
rect 21376 23032 21404 23063
rect 21545 23035 21603 23041
rect 21545 23032 21557 23035
rect 21376 23004 21557 23032
rect 20579 23001 20591 23004
rect 20533 22995 20591 23001
rect 21376 22976 21404 23004
rect 21545 23001 21557 23004
rect 21591 23001 21603 23035
rect 21545 22995 21603 23001
rect 21761 23035 21819 23041
rect 21761 23001 21773 23035
rect 21807 23032 21819 23035
rect 22066 23032 22094 23140
rect 22189 23137 22201 23140
rect 22235 23137 22247 23171
rect 22189 23131 22247 23137
rect 22296 23109 22324 23276
rect 22554 23264 22560 23316
rect 22612 23304 22618 23316
rect 22649 23307 22707 23313
rect 22649 23304 22661 23307
rect 22612 23276 22661 23304
rect 22612 23264 22618 23276
rect 22649 23273 22661 23276
rect 22695 23273 22707 23307
rect 22649 23267 22707 23273
rect 23109 23307 23167 23313
rect 23109 23273 23121 23307
rect 23155 23304 23167 23307
rect 23382 23304 23388 23316
rect 23155 23276 23388 23304
rect 23155 23273 23167 23276
rect 23109 23267 23167 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 23566 23264 23572 23316
rect 23624 23304 23630 23316
rect 23753 23307 23811 23313
rect 23753 23304 23765 23307
rect 23624 23276 23765 23304
rect 23624 23264 23630 23276
rect 23753 23273 23765 23276
rect 23799 23273 23811 23307
rect 23753 23267 23811 23273
rect 22370 23196 22376 23248
rect 22428 23236 22434 23248
rect 22428 23208 24072 23236
rect 22428 23196 22434 23208
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 22940 23140 23489 23168
rect 22940 23109 22968 23140
rect 23477 23137 23489 23140
rect 23523 23168 23535 23171
rect 23937 23171 23995 23177
rect 23937 23168 23949 23171
rect 23523 23140 23949 23168
rect 23523 23137 23535 23140
rect 23477 23131 23535 23137
rect 23937 23137 23949 23140
rect 23983 23137 23995 23171
rect 23937 23131 23995 23137
rect 22281 23103 22339 23109
rect 22281 23069 22293 23103
rect 22327 23100 22339 23103
rect 22925 23103 22983 23109
rect 22327 23072 22876 23100
rect 22327 23069 22339 23072
rect 22281 23063 22339 23069
rect 22554 23032 22560 23044
rect 21807 23004 22560 23032
rect 21807 23001 21819 23004
rect 21761 22995 21819 23001
rect 22554 22992 22560 23004
rect 22612 23032 22618 23044
rect 22741 23035 22799 23041
rect 22741 23032 22753 23035
rect 22612 23004 22753 23032
rect 22612 22992 22618 23004
rect 22741 23001 22753 23004
rect 22787 23001 22799 23035
rect 22848 23032 22876 23072
rect 22925 23069 22937 23103
rect 22971 23069 22983 23103
rect 22925 23063 22983 23069
rect 23385 23103 23443 23109
rect 23385 23069 23397 23103
rect 23431 23100 23443 23103
rect 23658 23100 23664 23112
rect 23431 23072 23664 23100
rect 23431 23069 23443 23072
rect 23385 23063 23443 23069
rect 23400 23032 23428 23063
rect 23658 23060 23664 23072
rect 23716 23060 23722 23112
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24044 23109 24072 23208
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23100 24087 23103
rect 24210 23100 24216 23112
rect 24075 23072 24216 23100
rect 24075 23069 24087 23072
rect 24029 23063 24087 23069
rect 24210 23060 24216 23072
rect 24268 23060 24274 23112
rect 22848 23004 23428 23032
rect 22741 22995 22799 23001
rect 17313 22967 17371 22973
rect 17313 22933 17325 22967
rect 17359 22933 17371 22967
rect 17313 22927 17371 22933
rect 17957 22967 18015 22973
rect 17957 22933 17969 22967
rect 18003 22964 18015 22967
rect 18230 22964 18236 22976
rect 18003 22936 18236 22964
rect 18003 22933 18015 22936
rect 17957 22927 18015 22933
rect 18230 22924 18236 22936
rect 18288 22924 18294 22976
rect 18322 22924 18328 22976
rect 18380 22924 18386 22976
rect 20898 22924 20904 22976
rect 20956 22964 20962 22976
rect 21358 22964 21364 22976
rect 20956 22936 21364 22964
rect 20956 22924 20962 22936
rect 21358 22924 21364 22936
rect 21416 22924 21422 22976
rect 1104 22874 26312 22896
rect 1104 22822 4761 22874
rect 4813 22822 4825 22874
rect 4877 22822 4889 22874
rect 4941 22822 4953 22874
rect 5005 22822 5017 22874
rect 5069 22822 11063 22874
rect 11115 22822 11127 22874
rect 11179 22822 11191 22874
rect 11243 22822 11255 22874
rect 11307 22822 11319 22874
rect 11371 22822 17365 22874
rect 17417 22822 17429 22874
rect 17481 22822 17493 22874
rect 17545 22822 17557 22874
rect 17609 22822 17621 22874
rect 17673 22822 23667 22874
rect 23719 22822 23731 22874
rect 23783 22822 23795 22874
rect 23847 22822 23859 22874
rect 23911 22822 23923 22874
rect 23975 22822 26312 22874
rect 1104 22800 26312 22822
rect 4062 22720 4068 22772
rect 4120 22720 4126 22772
rect 4985 22763 5043 22769
rect 4985 22729 4997 22763
rect 5031 22760 5043 22763
rect 6270 22760 6276 22772
rect 5031 22732 6276 22760
rect 5031 22729 5043 22732
rect 4985 22723 5043 22729
rect 6270 22720 6276 22732
rect 6328 22720 6334 22772
rect 9600 22732 9904 22760
rect 5994 22652 6000 22704
rect 6052 22692 6058 22704
rect 9214 22692 9220 22704
rect 6052 22664 9220 22692
rect 6052 22652 6058 22664
rect 9214 22652 9220 22664
rect 9272 22652 9278 22704
rect 9398 22652 9404 22704
rect 9456 22692 9462 22704
rect 9600 22701 9628 22732
rect 9585 22695 9643 22701
rect 9585 22692 9597 22695
rect 9456 22664 9597 22692
rect 9456 22652 9462 22664
rect 9585 22661 9597 22664
rect 9631 22661 9643 22695
rect 9585 22655 9643 22661
rect 9766 22652 9772 22704
rect 9824 22701 9830 22704
rect 9824 22695 9843 22701
rect 9831 22661 9843 22695
rect 9876 22692 9904 22732
rect 9950 22720 9956 22772
rect 10008 22720 10014 22772
rect 10778 22720 10784 22772
rect 10836 22760 10842 22772
rect 11165 22763 11223 22769
rect 11165 22760 11177 22763
rect 10836 22732 11177 22760
rect 10836 22720 10842 22732
rect 11165 22729 11177 22732
rect 11211 22729 11223 22763
rect 11165 22723 11223 22729
rect 11698 22720 11704 22772
rect 11756 22769 11762 22772
rect 11756 22763 11775 22769
rect 11763 22729 11775 22763
rect 11756 22723 11775 22729
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 11974 22760 11980 22772
rect 11931 22732 11980 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 11756 22720 11762 22723
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12066 22720 12072 22772
rect 12124 22760 12130 22772
rect 12453 22763 12511 22769
rect 12453 22760 12465 22763
rect 12124 22732 12465 22760
rect 12124 22720 12130 22732
rect 12453 22729 12465 22732
rect 12499 22729 12511 22763
rect 12453 22723 12511 22729
rect 12986 22720 12992 22772
rect 13044 22760 13050 22772
rect 13649 22763 13707 22769
rect 13649 22760 13661 22763
rect 13044 22732 13661 22760
rect 13044 22720 13050 22732
rect 13649 22729 13661 22732
rect 13695 22729 13707 22763
rect 13649 22723 13707 22729
rect 13817 22763 13875 22769
rect 13817 22729 13829 22763
rect 13863 22760 13875 22763
rect 13863 22732 18092 22760
rect 13863 22729 13875 22732
rect 13817 22723 13875 22729
rect 10965 22695 11023 22701
rect 10965 22692 10977 22695
rect 9876 22664 10977 22692
rect 9824 22655 9843 22661
rect 10965 22661 10977 22664
rect 11011 22661 11023 22695
rect 10965 22655 11023 22661
rect 11517 22695 11575 22701
rect 11517 22661 11529 22695
rect 11563 22661 11575 22695
rect 11517 22655 11575 22661
rect 12253 22695 12311 22701
rect 12253 22661 12265 22695
rect 12299 22692 12311 22695
rect 13449 22695 13507 22701
rect 13449 22692 13461 22695
rect 12299 22664 13461 22692
rect 12299 22661 12311 22664
rect 12253 22655 12311 22661
rect 13449 22661 13461 22664
rect 13495 22692 13507 22695
rect 15565 22695 15623 22701
rect 13495 22664 15424 22692
rect 13495 22661 13507 22664
rect 13449 22655 13507 22661
rect 9824 22652 9830 22655
rect 4249 22627 4307 22633
rect 4249 22593 4261 22627
rect 4295 22624 4307 22627
rect 4295 22596 4568 22624
rect 4295 22593 4307 22596
rect 4249 22587 4307 22593
rect 4540 22497 4568 22596
rect 4890 22584 4896 22636
rect 4948 22584 4954 22636
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22624 5779 22627
rect 6270 22624 6276 22636
rect 5767 22596 6276 22624
rect 5767 22593 5779 22596
rect 5721 22587 5779 22593
rect 6270 22584 6276 22596
rect 6328 22624 6334 22636
rect 6454 22624 6460 22636
rect 6328 22596 6460 22624
rect 6328 22584 6334 22596
rect 6454 22584 6460 22596
rect 6512 22584 6518 22636
rect 9232 22624 9260 22652
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 9232 22596 10241 22624
rect 10229 22593 10241 22596
rect 10275 22624 10287 22627
rect 10505 22627 10563 22633
rect 10505 22624 10517 22627
rect 10275 22596 10517 22624
rect 10275 22593 10287 22596
rect 10229 22587 10287 22593
rect 10505 22593 10517 22596
rect 10551 22593 10563 22627
rect 10980 22624 11008 22655
rect 11532 22624 11560 22655
rect 11606 22624 11612 22636
rect 10980 22596 11612 22624
rect 10505 22587 10563 22593
rect 11606 22584 11612 22596
rect 11664 22584 11670 22636
rect 11974 22584 11980 22636
rect 12032 22624 12038 22636
rect 12268 22624 12296 22655
rect 15010 22624 15016 22636
rect 12032 22596 12296 22624
rect 12636 22596 15016 22624
rect 12032 22584 12038 22596
rect 5169 22559 5227 22565
rect 5169 22525 5181 22559
rect 5215 22525 5227 22559
rect 12526 22556 12532 22568
rect 5169 22519 5227 22525
rect 12452 22528 12532 22556
rect 4525 22491 4583 22497
rect 4525 22457 4537 22491
rect 4571 22457 4583 22491
rect 5184 22488 5212 22519
rect 6178 22488 6184 22500
rect 5184 22460 6184 22488
rect 4525 22451 4583 22457
rect 6178 22448 6184 22460
rect 6236 22448 6242 22500
rect 12452 22488 12480 22528
rect 12526 22516 12532 22528
rect 12584 22516 12590 22568
rect 12636 22497 12664 22596
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 15396 22624 15424 22664
rect 15565 22661 15577 22695
rect 15611 22692 15623 22695
rect 15654 22692 15660 22704
rect 15611 22664 15660 22692
rect 15611 22661 15623 22664
rect 15565 22655 15623 22661
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 16209 22695 16267 22701
rect 16209 22661 16221 22695
rect 16255 22692 16267 22695
rect 16298 22692 16304 22704
rect 16255 22664 16304 22692
rect 16255 22661 16267 22664
rect 16209 22655 16267 22661
rect 16298 22652 16304 22664
rect 16356 22652 16362 22704
rect 17034 22652 17040 22704
rect 17092 22652 17098 22704
rect 15841 22627 15899 22633
rect 15841 22624 15853 22627
rect 15396 22596 15853 22624
rect 15841 22593 15853 22596
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 12802 22516 12808 22568
rect 12860 22556 12866 22568
rect 12986 22556 12992 22568
rect 12860 22528 12992 22556
rect 12860 22516 12866 22528
rect 12986 22516 12992 22528
rect 13044 22516 13050 22568
rect 15856 22556 15884 22587
rect 16390 22584 16396 22636
rect 16448 22624 16454 22636
rect 18064 22633 18092 22732
rect 18138 22720 18144 22772
rect 18196 22760 18202 22772
rect 18325 22763 18383 22769
rect 18325 22760 18337 22763
rect 18196 22732 18337 22760
rect 18196 22720 18202 22732
rect 18325 22729 18337 22732
rect 18371 22729 18383 22763
rect 18325 22723 18383 22729
rect 19702 22720 19708 22772
rect 19760 22720 19766 22772
rect 20070 22720 20076 22772
rect 20128 22760 20134 22772
rect 21450 22760 21456 22772
rect 20128 22732 21456 22760
rect 20128 22720 20134 22732
rect 21450 22720 21456 22732
rect 21508 22720 21514 22772
rect 22554 22720 22560 22772
rect 22612 22720 22618 22772
rect 18598 22652 18604 22704
rect 18656 22692 18662 22704
rect 18877 22695 18935 22701
rect 18877 22692 18889 22695
rect 18656 22664 18889 22692
rect 18656 22652 18662 22664
rect 18877 22661 18889 22664
rect 18923 22661 18935 22695
rect 19794 22692 19800 22704
rect 18877 22655 18935 22661
rect 19398 22664 19800 22692
rect 17405 22627 17463 22633
rect 17405 22624 17417 22627
rect 16448 22596 17417 22624
rect 16448 22584 16454 22596
rect 17405 22593 17417 22596
rect 17451 22593 17463 22627
rect 17405 22587 17463 22593
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22624 18199 22627
rect 18322 22624 18328 22636
rect 18187 22596 18328 22624
rect 18187 22593 18199 22596
rect 18141 22587 18199 22593
rect 16669 22559 16727 22565
rect 16669 22556 16681 22559
rect 15856 22528 16681 22556
rect 16669 22525 16681 22528
rect 16715 22556 16727 22559
rect 17126 22556 17132 22568
rect 16715 22528 17132 22556
rect 16715 22525 16727 22528
rect 16669 22519 16727 22525
rect 17126 22516 17132 22528
rect 17184 22556 17190 22568
rect 17310 22556 17316 22568
rect 17184 22528 17316 22556
rect 17184 22516 17190 22528
rect 17310 22516 17316 22528
rect 17368 22516 17374 22568
rect 17420 22556 17448 22587
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22624 18475 22627
rect 18506 22624 18512 22636
rect 18463 22596 18512 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19398 22633 19426 22664
rect 19794 22652 19800 22664
rect 19852 22652 19858 22704
rect 21542 22692 21548 22704
rect 21206 22664 21548 22692
rect 21542 22652 21548 22664
rect 21600 22652 21606 22704
rect 23750 22652 23756 22704
rect 23808 22652 23814 22704
rect 24210 22652 24216 22704
rect 24268 22692 24274 22704
rect 24443 22695 24501 22701
rect 24443 22692 24455 22695
rect 24268 22664 24455 22692
rect 24268 22652 24274 22664
rect 24443 22661 24455 22664
rect 24489 22661 24501 22695
rect 24443 22655 24501 22661
rect 19383 22627 19441 22633
rect 19383 22593 19395 22627
rect 19429 22593 19441 22627
rect 19383 22587 19441 22593
rect 19702 22584 19708 22636
rect 19760 22584 19766 22636
rect 22373 22627 22431 22633
rect 22373 22593 22385 22627
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 17957 22559 18015 22565
rect 17420 22528 17908 22556
rect 9784 22460 12480 22488
rect 12621 22491 12679 22497
rect 9784 22432 9812 22460
rect 9766 22380 9772 22432
rect 9824 22380 9830 22432
rect 10318 22380 10324 22432
rect 10376 22380 10382 22432
rect 10597 22423 10655 22429
rect 10597 22389 10609 22423
rect 10643 22420 10655 22423
rect 10870 22420 10876 22432
rect 10643 22392 10876 22420
rect 10643 22389 10655 22392
rect 10597 22383 10655 22389
rect 10870 22380 10876 22392
rect 10928 22380 10934 22432
rect 11164 22429 11192 22460
rect 11149 22423 11207 22429
rect 11149 22389 11161 22423
rect 11195 22389 11207 22423
rect 11149 22383 11207 22389
rect 11330 22380 11336 22432
rect 11388 22380 11394 22432
rect 11716 22429 11744 22460
rect 12621 22457 12633 22491
rect 12667 22457 12679 22491
rect 12621 22451 12679 22457
rect 12728 22460 13676 22488
rect 11701 22423 11759 22429
rect 11701 22389 11713 22423
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12728 22420 12756 22460
rect 12492 22392 12756 22420
rect 12492 22380 12498 22392
rect 12802 22380 12808 22432
rect 12860 22420 12866 22432
rect 13648 22429 13676 22460
rect 15194 22448 15200 22500
rect 15252 22448 15258 22500
rect 16022 22448 16028 22500
rect 16080 22488 16086 22500
rect 16393 22491 16451 22497
rect 16393 22488 16405 22491
rect 16080 22460 16405 22488
rect 16080 22448 16086 22460
rect 16393 22457 16405 22460
rect 16439 22457 16451 22491
rect 16393 22451 16451 22457
rect 17497 22491 17555 22497
rect 17497 22457 17509 22491
rect 17543 22488 17555 22491
rect 17770 22488 17776 22500
rect 17543 22460 17776 22488
rect 17543 22457 17555 22460
rect 17497 22451 17555 22457
rect 17770 22448 17776 22460
rect 17828 22448 17834 22500
rect 17880 22488 17908 22528
rect 17957 22525 17969 22559
rect 18003 22556 18015 22559
rect 19610 22556 19616 22568
rect 18003 22528 19104 22556
rect 18003 22525 18015 22528
rect 17957 22519 18015 22525
rect 18322 22488 18328 22500
rect 17880 22460 18328 22488
rect 18322 22448 18328 22460
rect 18380 22488 18386 22500
rect 19076 22497 19104 22528
rect 19444 22528 19616 22556
rect 19444 22500 19472 22528
rect 19610 22516 19616 22528
rect 19668 22556 19674 22568
rect 19797 22559 19855 22565
rect 19797 22556 19809 22559
rect 19668 22528 19809 22556
rect 19668 22516 19674 22528
rect 19797 22525 19809 22528
rect 19843 22525 19855 22559
rect 19797 22519 19855 22525
rect 20165 22559 20223 22565
rect 20165 22525 20177 22559
rect 20211 22556 20223 22559
rect 20346 22556 20352 22568
rect 20211 22528 20352 22556
rect 20211 22525 20223 22528
rect 20165 22519 20223 22525
rect 20346 22516 20352 22528
rect 20404 22516 20410 22568
rect 20990 22516 20996 22568
rect 21048 22556 21054 22568
rect 22189 22559 22247 22565
rect 22189 22556 22201 22559
rect 21048 22528 22201 22556
rect 21048 22516 21054 22528
rect 22189 22525 22201 22528
rect 22235 22556 22247 22559
rect 22278 22556 22284 22568
rect 22235 22528 22284 22556
rect 22235 22525 22247 22528
rect 22189 22519 22247 22525
rect 22278 22516 22284 22528
rect 22336 22516 22342 22568
rect 22388 22556 22416 22587
rect 22646 22584 22652 22636
rect 22704 22584 22710 22636
rect 22922 22584 22928 22636
rect 22980 22624 22986 22636
rect 23017 22627 23075 22633
rect 23017 22624 23029 22627
rect 22980 22596 23029 22624
rect 22980 22584 22986 22596
rect 23017 22593 23029 22596
rect 23063 22593 23075 22627
rect 23017 22587 23075 22593
rect 24026 22556 24032 22568
rect 22388 22528 24032 22556
rect 18509 22491 18567 22497
rect 18509 22488 18521 22491
rect 18380 22460 18521 22488
rect 18380 22448 18386 22460
rect 18509 22457 18521 22460
rect 18555 22457 18567 22491
rect 18509 22451 18567 22457
rect 19061 22491 19119 22497
rect 19061 22457 19073 22491
rect 19107 22457 19119 22491
rect 19061 22451 19119 22457
rect 19426 22448 19432 22500
rect 19484 22448 19490 22500
rect 21358 22448 21364 22500
rect 21416 22488 21422 22500
rect 21591 22491 21649 22497
rect 21591 22488 21603 22491
rect 21416 22460 21603 22488
rect 21416 22448 21422 22460
rect 21591 22457 21603 22460
rect 21637 22457 21649 22491
rect 21591 22451 21649 22457
rect 13357 22423 13415 22429
rect 13357 22420 13369 22423
rect 12860 22392 13369 22420
rect 12860 22380 12866 22392
rect 13357 22389 13369 22392
rect 13403 22389 13415 22423
rect 13357 22383 13415 22389
rect 13633 22423 13691 22429
rect 13633 22389 13645 22423
rect 13679 22420 13691 22423
rect 13722 22420 13728 22432
rect 13679 22392 13728 22420
rect 13679 22389 13691 22392
rect 13633 22383 13691 22389
rect 13722 22380 13728 22392
rect 13780 22380 13786 22432
rect 15562 22380 15568 22432
rect 15620 22380 15626 22432
rect 15749 22423 15807 22429
rect 15749 22389 15761 22423
rect 15795 22420 15807 22423
rect 16114 22420 16120 22432
rect 15795 22392 16120 22420
rect 15795 22389 15807 22392
rect 15749 22383 15807 22389
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16209 22423 16267 22429
rect 16209 22389 16221 22423
rect 16255 22420 16267 22423
rect 16298 22420 16304 22432
rect 16255 22392 16304 22420
rect 16255 22389 16267 22392
rect 16209 22383 16267 22389
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 17034 22380 17040 22432
rect 17092 22380 17098 22432
rect 17218 22380 17224 22432
rect 17276 22380 17282 22432
rect 17678 22380 17684 22432
rect 17736 22380 17742 22432
rect 18874 22380 18880 22432
rect 18932 22380 18938 22432
rect 19521 22423 19579 22429
rect 19521 22389 19533 22423
rect 19567 22420 19579 22423
rect 19702 22420 19708 22432
rect 19567 22392 19708 22420
rect 19567 22389 19579 22392
rect 19521 22383 19579 22389
rect 19702 22380 19708 22392
rect 19760 22420 19766 22432
rect 21082 22420 21088 22432
rect 19760 22392 21088 22420
rect 19760 22380 19766 22392
rect 21082 22380 21088 22392
rect 21140 22420 21146 22432
rect 22388 22420 22416 22528
rect 24026 22516 24032 22528
rect 24084 22516 24090 22568
rect 21140 22392 22416 22420
rect 21140 22380 21146 22392
rect 1104 22330 26312 22352
rect 1104 22278 4101 22330
rect 4153 22278 4165 22330
rect 4217 22278 4229 22330
rect 4281 22278 4293 22330
rect 4345 22278 4357 22330
rect 4409 22278 10403 22330
rect 10455 22278 10467 22330
rect 10519 22278 10531 22330
rect 10583 22278 10595 22330
rect 10647 22278 10659 22330
rect 10711 22278 16705 22330
rect 16757 22278 16769 22330
rect 16821 22278 16833 22330
rect 16885 22278 16897 22330
rect 16949 22278 16961 22330
rect 17013 22278 23007 22330
rect 23059 22278 23071 22330
rect 23123 22278 23135 22330
rect 23187 22278 23199 22330
rect 23251 22278 23263 22330
rect 23315 22278 26312 22330
rect 1104 22256 26312 22278
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 11388 22188 14964 22216
rect 11388 22176 11394 22188
rect 11149 22151 11207 22157
rect 11149 22117 11161 22151
rect 11195 22148 11207 22151
rect 11974 22148 11980 22160
rect 11195 22120 11980 22148
rect 11195 22117 11207 22120
rect 11149 22111 11207 22117
rect 11974 22108 11980 22120
rect 12032 22108 12038 22160
rect 14936 22148 14964 22188
rect 15930 22176 15936 22228
rect 15988 22176 15994 22228
rect 16485 22219 16543 22225
rect 16485 22185 16497 22219
rect 16531 22216 16543 22219
rect 17126 22216 17132 22228
rect 16531 22188 17132 22216
rect 16531 22185 16543 22188
rect 16485 22179 16543 22185
rect 17126 22176 17132 22188
rect 17184 22176 17190 22228
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 17589 22219 17647 22225
rect 17589 22216 17601 22219
rect 17276 22188 17601 22216
rect 17276 22176 17282 22188
rect 17589 22185 17601 22188
rect 17635 22185 17647 22219
rect 17589 22179 17647 22185
rect 17681 22219 17739 22225
rect 17681 22185 17693 22219
rect 17727 22216 17739 22219
rect 17862 22216 17868 22228
rect 17727 22188 17868 22216
rect 17727 22185 17739 22188
rect 17681 22179 17739 22185
rect 17862 22176 17868 22188
rect 17920 22176 17926 22228
rect 18064 22188 18460 22216
rect 17497 22151 17555 22157
rect 17497 22148 17509 22151
rect 14936 22120 17509 22148
rect 17497 22117 17509 22120
rect 17543 22117 17555 22151
rect 17497 22111 17555 22117
rect 17770 22108 17776 22160
rect 17828 22148 17834 22160
rect 18064 22148 18092 22188
rect 17828 22120 18092 22148
rect 17828 22108 17834 22120
rect 18322 22108 18328 22160
rect 18380 22108 18386 22160
rect 18432 22148 18460 22188
rect 18506 22176 18512 22228
rect 18564 22176 18570 22228
rect 18785 22219 18843 22225
rect 18785 22185 18797 22219
rect 18831 22185 18843 22219
rect 18785 22179 18843 22185
rect 18800 22148 18828 22179
rect 19242 22176 19248 22228
rect 19300 22216 19306 22228
rect 19705 22219 19763 22225
rect 19705 22216 19717 22219
rect 19300 22188 19717 22216
rect 19300 22176 19306 22188
rect 19705 22185 19717 22188
rect 19751 22185 19763 22219
rect 19705 22179 19763 22185
rect 20070 22176 20076 22228
rect 20128 22216 20134 22228
rect 20165 22219 20223 22225
rect 20165 22216 20177 22219
rect 20128 22188 20177 22216
rect 20128 22176 20134 22188
rect 20165 22185 20177 22188
rect 20211 22185 20223 22219
rect 20165 22179 20223 22185
rect 18432 22120 18828 22148
rect 5813 22083 5871 22089
rect 5813 22049 5825 22083
rect 5859 22080 5871 22083
rect 12710 22080 12716 22092
rect 5859 22052 6040 22080
rect 5859 22049 5871 22052
rect 5813 22043 5871 22049
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 22012 3847 22015
rect 4154 22012 4160 22024
rect 3835 21984 4160 22012
rect 3835 21981 3847 21984
rect 3789 21975 3847 21981
rect 4154 21972 4160 21984
rect 4212 21972 4218 22024
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 5902 21972 5908 22024
rect 5960 21972 5966 22024
rect 6012 22021 6040 22052
rect 11440 22052 12716 22080
rect 5997 22015 6055 22021
rect 5997 21981 6009 22015
rect 6043 21981 6055 22015
rect 5997 21975 6055 21981
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6181 21975 6239 21981
rect 6196 21944 6224 21975
rect 6730 21972 6736 22024
rect 6788 22012 6794 22024
rect 6917 22015 6975 22021
rect 6917 22012 6929 22015
rect 6788 21984 6929 22012
rect 6788 21972 6794 21984
rect 6917 21981 6929 21984
rect 6963 21981 6975 22015
rect 6917 21975 6975 21981
rect 8754 21972 8760 22024
rect 8812 21972 8818 22024
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 9306 21972 9312 22024
rect 9364 22012 9370 22024
rect 11440 22021 11468 22052
rect 12710 22040 12716 22052
rect 12768 22040 12774 22092
rect 12986 22040 12992 22092
rect 13044 22080 13050 22092
rect 13817 22083 13875 22089
rect 13817 22080 13829 22083
rect 13044 22052 13829 22080
rect 13044 22040 13050 22052
rect 13817 22049 13829 22052
rect 13863 22049 13875 22083
rect 13817 22043 13875 22049
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 9364 21984 9413 22012
rect 9364 21972 9370 21984
rect 9401 21981 9413 21984
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 11425 22015 11483 22021
rect 11425 21981 11437 22015
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 11701 22015 11759 22021
rect 11701 21981 11713 22015
rect 11747 22012 11759 22015
rect 11974 22012 11980 22024
rect 11747 21984 11980 22012
rect 11747 21981 11759 21984
rect 11701 21975 11759 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 7466 21944 7472 21956
rect 6196 21916 7472 21944
rect 7466 21904 7472 21916
rect 7524 21904 7530 21956
rect 9677 21947 9735 21953
rect 9677 21944 9689 21947
rect 8588 21916 9689 21944
rect 3786 21836 3792 21888
rect 3844 21876 3850 21888
rect 3973 21879 4031 21885
rect 3973 21876 3985 21879
rect 3844 21848 3985 21876
rect 3844 21836 3850 21848
rect 3973 21845 3985 21848
rect 4019 21845 4031 21879
rect 3973 21839 4031 21845
rect 6181 21879 6239 21885
rect 6181 21845 6193 21879
rect 6227 21876 6239 21879
rect 6638 21876 6644 21888
rect 6227 21848 6644 21876
rect 6227 21845 6239 21848
rect 6181 21839 6239 21845
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 7009 21879 7067 21885
rect 7009 21845 7021 21879
rect 7055 21876 7067 21879
rect 7098 21876 7104 21888
rect 7055 21848 7104 21876
rect 7055 21845 7067 21848
rect 7009 21839 7067 21845
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 8588 21885 8616 21916
rect 9677 21913 9689 21916
rect 9723 21913 9735 21947
rect 9677 21907 9735 21913
rect 10318 21904 10324 21956
rect 10376 21904 10382 21956
rect 11517 21947 11575 21953
rect 11517 21913 11529 21947
rect 11563 21944 11575 21947
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 11563 21916 12357 21944
rect 11563 21913 11575 21916
rect 11517 21907 11575 21913
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 12345 21907 12403 21913
rect 13078 21904 13084 21956
rect 13136 21904 13142 21956
rect 13832 21944 13860 22043
rect 15010 22040 15016 22092
rect 15068 22080 15074 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15068 22052 15761 22080
rect 15068 22040 15074 22052
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 15749 22043 15807 22049
rect 16114 22040 16120 22092
rect 16172 22080 16178 22092
rect 16301 22083 16359 22089
rect 16301 22080 16313 22083
rect 16172 22052 16313 22080
rect 16172 22040 16178 22052
rect 16301 22049 16313 22052
rect 16347 22049 16359 22083
rect 17310 22080 17316 22092
rect 16301 22043 16359 22049
rect 17052 22052 17316 22080
rect 13906 21972 13912 22024
rect 13964 22012 13970 22024
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13964 21984 14105 22012
rect 13964 21972 13970 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14274 21972 14280 22024
rect 14332 22012 14338 22024
rect 14461 22015 14519 22021
rect 14461 22012 14473 22015
rect 14332 21984 14473 22012
rect 14332 21972 14338 21984
rect 14461 21981 14473 21984
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 15197 22015 15255 22021
rect 15197 22012 15209 22015
rect 15151 21984 15209 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 15197 21981 15209 21984
rect 15243 21981 15255 22015
rect 15197 21975 15255 21981
rect 15286 21972 15292 22024
rect 15344 21972 15350 22024
rect 15933 22015 15991 22021
rect 15933 21981 15945 22015
rect 15979 22012 15991 22015
rect 15979 21984 16160 22012
rect 15979 21981 15991 21984
rect 15933 21975 15991 21981
rect 15304 21944 15332 21972
rect 13832 21916 15332 21944
rect 15657 21947 15715 21953
rect 15657 21913 15669 21947
rect 15703 21944 15715 21947
rect 16022 21944 16028 21956
rect 15703 21916 16028 21944
rect 15703 21913 15715 21916
rect 15657 21907 15715 21913
rect 16022 21904 16028 21916
rect 16080 21904 16086 21956
rect 16132 21944 16160 21984
rect 16206 21972 16212 22024
rect 16264 21972 16270 22024
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 16500 21944 16528 21975
rect 16850 21972 16856 22024
rect 16908 21972 16914 22024
rect 17052 22021 17080 22052
rect 17310 22040 17316 22052
rect 17368 22080 17374 22092
rect 18049 22083 18107 22089
rect 18049 22080 18061 22083
rect 17368 22052 18061 22080
rect 17368 22040 17374 22052
rect 18049 22049 18061 22052
rect 18095 22049 18107 22083
rect 18049 22043 18107 22049
rect 19794 22040 19800 22092
rect 19852 22040 19858 22092
rect 21542 22040 21548 22092
rect 21600 22040 21606 22092
rect 23750 22040 23756 22092
rect 23808 22040 23814 22092
rect 17037 22015 17095 22021
rect 17037 21981 17049 22015
rect 17083 21981 17095 22015
rect 17037 21975 17095 21981
rect 17770 21972 17776 22024
rect 17828 21972 17834 22024
rect 17957 22015 18015 22021
rect 17957 21981 17969 22015
rect 18003 22012 18015 22015
rect 19242 22012 19248 22024
rect 18003 21984 19248 22012
rect 18003 21981 18015 21984
rect 17957 21975 18015 21981
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19518 21972 19524 22024
rect 19576 22012 19582 22024
rect 19981 22015 20039 22021
rect 19981 22012 19993 22015
rect 19576 21984 19993 22012
rect 19576 21972 19582 21984
rect 19981 21981 19993 21984
rect 20027 21981 20039 22015
rect 19981 21975 20039 21981
rect 21453 22015 21511 22021
rect 21453 21981 21465 22015
rect 21499 22012 21511 22015
rect 23661 22015 23719 22021
rect 23661 22012 23673 22015
rect 21499 21984 23673 22012
rect 21499 21981 21511 21984
rect 21453 21975 21511 21981
rect 23661 21981 23673 21984
rect 23707 22012 23719 22015
rect 24302 22012 24308 22024
rect 23707 21984 24308 22012
rect 23707 21981 23719 21984
rect 23661 21975 23719 21981
rect 24302 21972 24308 21984
rect 24360 21972 24366 22024
rect 16945 21947 17003 21953
rect 16945 21944 16957 21947
rect 16132 21916 16957 21944
rect 16945 21913 16957 21916
rect 16991 21944 17003 21947
rect 17862 21944 17868 21956
rect 16991 21916 17868 21944
rect 16991 21913 17003 21916
rect 16945 21907 17003 21913
rect 17862 21904 17868 21916
rect 17920 21904 17926 21956
rect 18046 21904 18052 21956
rect 18104 21944 18110 21956
rect 18598 21944 18604 21956
rect 18104 21916 18604 21944
rect 18104 21904 18110 21916
rect 18598 21904 18604 21916
rect 18656 21904 18662 21956
rect 18817 21947 18875 21953
rect 18817 21913 18829 21947
rect 18863 21944 18875 21947
rect 18863 21916 19656 21944
rect 18863 21913 18875 21916
rect 18817 21907 18875 21913
rect 8573 21879 8631 21885
rect 8573 21845 8585 21879
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 8938 21836 8944 21888
rect 8996 21836 9002 21888
rect 11606 21836 11612 21888
rect 11664 21876 11670 21888
rect 11885 21879 11943 21885
rect 11885 21876 11897 21879
rect 11664 21848 11897 21876
rect 11664 21836 11670 21848
rect 11885 21845 11897 21848
rect 11931 21845 11943 21879
rect 11885 21839 11943 21845
rect 12526 21836 12532 21888
rect 12584 21876 12590 21888
rect 13630 21876 13636 21888
rect 12584 21848 13636 21876
rect 12584 21836 12590 21848
rect 13630 21836 13636 21848
rect 13688 21876 13694 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13688 21848 14289 21876
rect 13688 21836 13694 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 14277 21839 14335 21845
rect 14458 21836 14464 21888
rect 14516 21876 14522 21888
rect 15289 21879 15347 21885
rect 15289 21876 15301 21879
rect 14516 21848 15301 21876
rect 14516 21836 14522 21848
rect 15289 21845 15301 21848
rect 15335 21845 15347 21879
rect 15289 21839 15347 21845
rect 16117 21879 16175 21885
rect 16117 21845 16129 21879
rect 16163 21876 16175 21879
rect 16206 21876 16212 21888
rect 16163 21848 16212 21876
rect 16163 21845 16175 21848
rect 16117 21839 16175 21845
rect 16206 21836 16212 21848
rect 16264 21836 16270 21888
rect 16574 21836 16580 21888
rect 16632 21876 16638 21888
rect 16669 21879 16727 21885
rect 16669 21876 16681 21879
rect 16632 21848 16681 21876
rect 16632 21836 16638 21848
rect 16669 21845 16681 21848
rect 16715 21845 16727 21879
rect 16669 21839 16727 21845
rect 17034 21836 17040 21888
rect 17092 21876 17098 21888
rect 17221 21879 17279 21885
rect 17221 21876 17233 21879
rect 17092 21848 17233 21876
rect 17092 21836 17098 21848
rect 17221 21845 17233 21848
rect 17267 21845 17279 21879
rect 17221 21839 17279 21845
rect 18966 21836 18972 21888
rect 19024 21836 19030 21888
rect 19628 21876 19656 21916
rect 19702 21904 19708 21956
rect 19760 21904 19766 21956
rect 21082 21876 21088 21888
rect 19628 21848 21088 21876
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 1104 21786 26312 21808
rect 1104 21734 4761 21786
rect 4813 21734 4825 21786
rect 4877 21734 4889 21786
rect 4941 21734 4953 21786
rect 5005 21734 5017 21786
rect 5069 21734 11063 21786
rect 11115 21734 11127 21786
rect 11179 21734 11191 21786
rect 11243 21734 11255 21786
rect 11307 21734 11319 21786
rect 11371 21734 17365 21786
rect 17417 21734 17429 21786
rect 17481 21734 17493 21786
rect 17545 21734 17557 21786
rect 17609 21734 17621 21786
rect 17673 21734 23667 21786
rect 23719 21734 23731 21786
rect 23783 21734 23795 21786
rect 23847 21734 23859 21786
rect 23911 21734 23923 21786
rect 23975 21734 26312 21786
rect 1104 21712 26312 21734
rect 3602 21632 3608 21684
rect 3660 21672 3666 21684
rect 5534 21672 5540 21684
rect 3660 21644 5540 21672
rect 3660 21632 3666 21644
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 8389 21675 8447 21681
rect 8389 21641 8401 21675
rect 8435 21672 8447 21675
rect 9122 21672 9128 21684
rect 8435 21644 9128 21672
rect 8435 21641 8447 21644
rect 8389 21635 8447 21641
rect 9122 21632 9128 21644
rect 9180 21632 9186 21684
rect 12434 21672 12440 21684
rect 11348 21644 12440 21672
rect 2498 21564 2504 21616
rect 2556 21564 2562 21616
rect 3510 21564 3516 21616
rect 3568 21604 3574 21616
rect 3568 21576 4370 21604
rect 3568 21564 3574 21576
rect 6638 21564 6644 21616
rect 6696 21564 6702 21616
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 8938 21564 8944 21616
rect 8996 21604 9002 21616
rect 9585 21607 9643 21613
rect 9585 21604 9597 21607
rect 8996 21576 9597 21604
rect 8996 21564 9002 21576
rect 9585 21573 9597 21576
rect 9631 21573 9643 21607
rect 10870 21604 10876 21616
rect 10810 21576 10876 21604
rect 9585 21567 9643 21573
rect 10870 21564 10876 21576
rect 10928 21564 10934 21616
rect 11348 21613 11376 21644
rect 12434 21632 12440 21644
rect 12492 21632 12498 21684
rect 13722 21632 13728 21684
rect 13780 21672 13786 21684
rect 16298 21672 16304 21684
rect 13780 21644 16304 21672
rect 13780 21632 13786 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 17126 21632 17132 21684
rect 17184 21672 17190 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 17184 21644 17693 21672
rect 17184 21632 17190 21644
rect 17681 21641 17693 21644
rect 17727 21641 17739 21675
rect 17681 21635 17739 21641
rect 11333 21607 11391 21613
rect 11333 21573 11345 21607
rect 11379 21573 11391 21607
rect 14366 21604 14372 21616
rect 13846 21576 14372 21604
rect 11333 21567 11391 21573
rect 14366 21564 14372 21576
rect 14424 21564 14430 21616
rect 16114 21564 16120 21616
rect 16172 21604 16178 21616
rect 17497 21607 17555 21613
rect 17497 21604 17509 21607
rect 16172 21576 17509 21604
rect 16172 21564 16178 21576
rect 17497 21573 17509 21576
rect 17543 21604 17555 21607
rect 18046 21604 18052 21616
rect 17543 21576 18052 21604
rect 17543 21573 17555 21576
rect 17497 21567 17555 21573
rect 18046 21564 18052 21576
rect 18104 21564 18110 21616
rect 18966 21604 18972 21616
rect 18156 21576 18972 21604
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 8662 21496 8668 21548
rect 8720 21536 8726 21548
rect 8757 21539 8815 21545
rect 8757 21536 8769 21539
rect 8720 21508 8769 21536
rect 8720 21496 8726 21508
rect 8757 21505 8769 21508
rect 8803 21505 8815 21539
rect 8757 21499 8815 21505
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21536 8907 21539
rect 8895 21508 9260 21536
rect 8895 21505 8907 21508
rect 8849 21499 8907 21505
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 1489 21471 1547 21477
rect 1489 21468 1501 21471
rect 1452 21440 1501 21468
rect 1452 21428 1458 21440
rect 1489 21437 1501 21440
rect 1535 21437 1547 21471
rect 1489 21431 1547 21437
rect 1765 21471 1823 21477
rect 1765 21437 1777 21471
rect 1811 21468 1823 21471
rect 2130 21468 2136 21480
rect 1811 21440 2136 21468
rect 1811 21437 1823 21440
rect 1765 21431 1823 21437
rect 1504 21332 1532 21431
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 3513 21471 3571 21477
rect 3513 21437 3525 21471
rect 3559 21437 3571 21471
rect 3513 21431 3571 21437
rect 2866 21360 2872 21412
rect 2924 21400 2930 21412
rect 3528 21400 3556 21431
rect 3878 21428 3884 21480
rect 3936 21428 3942 21480
rect 5166 21428 5172 21480
rect 5224 21468 5230 21480
rect 5353 21471 5411 21477
rect 5353 21468 5365 21471
rect 5224 21440 5365 21468
rect 5224 21428 5230 21440
rect 5353 21437 5365 21440
rect 5399 21468 5411 21471
rect 5537 21471 5595 21477
rect 5537 21468 5549 21471
rect 5399 21440 5549 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 5537 21437 5549 21440
rect 5583 21437 5595 21471
rect 5537 21431 5595 21437
rect 5626 21428 5632 21480
rect 5684 21468 5690 21480
rect 6362 21468 6368 21480
rect 5684 21440 6368 21468
rect 5684 21428 5690 21440
rect 6362 21428 6368 21440
rect 6420 21428 6426 21480
rect 8941 21471 8999 21477
rect 8941 21437 8953 21471
rect 8987 21437 8999 21471
rect 8941 21431 8999 21437
rect 6181 21403 6239 21409
rect 6181 21400 6193 21403
rect 2924 21372 3556 21400
rect 4908 21372 6193 21400
rect 2924 21360 2930 21372
rect 3602 21332 3608 21344
rect 1504 21304 3608 21332
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 3970 21292 3976 21344
rect 4028 21332 4034 21344
rect 4908 21332 4936 21372
rect 6181 21369 6193 21372
rect 6227 21369 6239 21403
rect 6181 21363 6239 21369
rect 8018 21360 8024 21412
rect 8076 21400 8082 21412
rect 8956 21400 8984 21431
rect 8076 21372 8984 21400
rect 8076 21360 8082 21372
rect 4028 21304 4936 21332
rect 4028 21292 4034 21304
rect 7650 21292 7656 21344
rect 7708 21332 7714 21344
rect 8113 21335 8171 21341
rect 8113 21332 8125 21335
rect 7708 21304 8125 21332
rect 7708 21292 7714 21304
rect 8113 21301 8125 21304
rect 8159 21301 8171 21335
rect 9232 21332 9260 21508
rect 12066 21496 12072 21548
rect 12124 21536 12130 21548
rect 12437 21539 12495 21545
rect 12437 21536 12449 21539
rect 12124 21508 12449 21536
rect 12124 21496 12130 21508
rect 12437 21505 12449 21508
rect 12483 21505 12495 21539
rect 14458 21536 14464 21548
rect 12437 21499 12495 21505
rect 14016 21508 14464 21536
rect 9306 21428 9312 21480
rect 9364 21428 9370 21480
rect 12805 21471 12863 21477
rect 12805 21437 12817 21471
rect 12851 21468 12863 21471
rect 14016 21468 14044 21508
rect 14458 21496 14464 21508
rect 14516 21496 14522 21548
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 14734 21536 14740 21548
rect 14599 21508 14740 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 15286 21496 15292 21548
rect 15344 21496 15350 21548
rect 15562 21496 15568 21548
rect 15620 21496 15626 21548
rect 18156 21545 18184 21576
rect 18966 21564 18972 21576
rect 19024 21564 19030 21616
rect 18141 21539 18199 21545
rect 18141 21505 18153 21539
rect 18187 21505 18199 21539
rect 18141 21499 18199 21505
rect 18230 21496 18236 21548
rect 18288 21536 18294 21548
rect 18325 21539 18383 21545
rect 18325 21536 18337 21539
rect 18288 21508 18337 21536
rect 18288 21496 18294 21508
rect 18325 21505 18337 21508
rect 18371 21505 18383 21539
rect 18325 21499 18383 21505
rect 18598 21496 18604 21548
rect 18656 21496 18662 21548
rect 25774 21496 25780 21548
rect 25832 21496 25838 21548
rect 12851 21440 14044 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 14090 21428 14096 21480
rect 14148 21468 14154 21480
rect 14369 21471 14427 21477
rect 14369 21468 14381 21471
rect 14148 21440 14381 21468
rect 14148 21428 14154 21440
rect 14369 21437 14381 21440
rect 14415 21437 14427 21471
rect 15406 21471 15464 21477
rect 15406 21468 15418 21471
rect 14369 21431 14427 21437
rect 14936 21440 15418 21468
rect 14274 21409 14280 21412
rect 14231 21403 14280 21409
rect 14231 21369 14243 21403
rect 14277 21369 14280 21403
rect 14231 21363 14280 21369
rect 14274 21360 14280 21363
rect 14332 21400 14338 21412
rect 14936 21400 14964 21440
rect 15406 21437 15418 21440
rect 15452 21437 15464 21471
rect 15580 21468 15608 21496
rect 16850 21468 16856 21480
rect 15580 21440 16856 21468
rect 15406 21431 15464 21437
rect 16850 21428 16856 21440
rect 16908 21468 16914 21480
rect 17129 21471 17187 21477
rect 17129 21468 17141 21471
rect 16908 21440 17141 21468
rect 16908 21428 16914 21440
rect 17129 21437 17141 21440
rect 17175 21468 17187 21471
rect 17494 21468 17500 21480
rect 17175 21440 17500 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 17494 21428 17500 21440
rect 17552 21428 17558 21480
rect 18417 21471 18475 21477
rect 18417 21437 18429 21471
rect 18463 21468 18475 21471
rect 19978 21468 19984 21480
rect 18463 21440 19984 21468
rect 18463 21437 18475 21440
rect 18417 21431 18475 21437
rect 19978 21428 19984 21440
rect 20036 21468 20042 21480
rect 21358 21468 21364 21480
rect 20036 21440 21364 21468
rect 20036 21428 20042 21440
rect 21358 21428 21364 21440
rect 21416 21428 21422 21480
rect 14332 21372 14964 21400
rect 15013 21403 15071 21409
rect 14332 21360 14338 21372
rect 15013 21369 15025 21403
rect 15059 21400 15071 21403
rect 15102 21400 15108 21412
rect 15059 21372 15108 21400
rect 15059 21369 15071 21372
rect 15013 21363 15071 21369
rect 15102 21360 15108 21372
rect 15160 21360 15166 21412
rect 17512 21372 18092 21400
rect 9766 21332 9772 21344
rect 9232 21304 9772 21332
rect 8113 21295 8171 21301
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 13630 21292 13636 21344
rect 13688 21332 13694 21344
rect 15562 21332 15568 21344
rect 13688 21304 15568 21332
rect 13688 21292 13694 21304
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 17512 21341 17540 21372
rect 16209 21335 16267 21341
rect 16209 21332 16221 21335
rect 16080 21304 16221 21332
rect 16080 21292 16086 21304
rect 16209 21301 16221 21304
rect 16255 21301 16267 21335
rect 16209 21295 16267 21301
rect 17497 21335 17555 21341
rect 17497 21301 17509 21335
rect 17543 21301 17555 21335
rect 17497 21295 17555 21301
rect 17862 21292 17868 21344
rect 17920 21332 17926 21344
rect 17957 21335 18015 21341
rect 17957 21332 17969 21335
rect 17920 21304 17969 21332
rect 17920 21292 17926 21304
rect 17957 21301 17969 21304
rect 18003 21301 18015 21335
rect 18064 21332 18092 21372
rect 18138 21360 18144 21412
rect 18196 21400 18202 21412
rect 18233 21403 18291 21409
rect 18233 21400 18245 21403
rect 18196 21372 18245 21400
rect 18196 21360 18202 21372
rect 18233 21369 18245 21372
rect 18279 21369 18291 21403
rect 18233 21363 18291 21369
rect 19794 21332 19800 21344
rect 18064 21304 19800 21332
rect 17957 21295 18015 21301
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 25958 21292 25964 21344
rect 26016 21292 26022 21344
rect 1104 21242 26312 21264
rect 1104 21190 4101 21242
rect 4153 21190 4165 21242
rect 4217 21190 4229 21242
rect 4281 21190 4293 21242
rect 4345 21190 4357 21242
rect 4409 21190 10403 21242
rect 10455 21190 10467 21242
rect 10519 21190 10531 21242
rect 10583 21190 10595 21242
rect 10647 21190 10659 21242
rect 10711 21190 16705 21242
rect 16757 21190 16769 21242
rect 16821 21190 16833 21242
rect 16885 21190 16897 21242
rect 16949 21190 16961 21242
rect 17013 21190 23007 21242
rect 23059 21190 23071 21242
rect 23123 21190 23135 21242
rect 23187 21190 23199 21242
rect 23251 21190 23263 21242
rect 23315 21190 26312 21242
rect 1104 21168 26312 21190
rect 2130 21088 2136 21140
rect 2188 21088 2194 21140
rect 2498 21088 2504 21140
rect 2556 21088 2562 21140
rect 2774 21128 2780 21140
rect 2700 21100 2780 21128
rect 1949 20995 2007 21001
rect 1949 20961 1961 20995
rect 1995 20992 2007 20995
rect 2700 20992 2728 21100
rect 2774 21088 2780 21100
rect 2832 21128 2838 21140
rect 3418 21128 3424 21140
rect 2832 21100 3424 21128
rect 2832 21088 2838 21100
rect 3418 21088 3424 21100
rect 3476 21088 3482 21140
rect 3510 21088 3516 21140
rect 3568 21088 3574 21140
rect 3789 21131 3847 21137
rect 3789 21097 3801 21131
rect 3835 21128 3847 21131
rect 3878 21128 3884 21140
rect 3835 21100 3884 21128
rect 3835 21097 3847 21100
rect 3789 21091 3847 21097
rect 3878 21088 3884 21100
rect 3936 21088 3942 21140
rect 4338 21088 4344 21140
rect 4396 21128 4402 21140
rect 4893 21131 4951 21137
rect 4893 21128 4905 21131
rect 4396 21100 4905 21128
rect 4396 21088 4402 21100
rect 4893 21097 4905 21100
rect 4939 21097 4951 21131
rect 4893 21091 4951 21097
rect 5077 21131 5135 21137
rect 5077 21097 5089 21131
rect 5123 21128 5135 21131
rect 5258 21128 5264 21140
rect 5123 21100 5264 21128
rect 5123 21097 5135 21100
rect 5077 21091 5135 21097
rect 5258 21088 5264 21100
rect 5316 21128 5322 21140
rect 5626 21128 5632 21140
rect 5316 21100 5632 21128
rect 5316 21088 5322 21100
rect 5626 21088 5632 21100
rect 5684 21088 5690 21140
rect 5902 21128 5908 21140
rect 5736 21100 5908 21128
rect 4525 21063 4583 21069
rect 4525 21029 4537 21063
rect 4571 21060 4583 21063
rect 5166 21060 5172 21072
rect 4571 21032 5172 21060
rect 4571 21029 4583 21032
rect 4525 21023 4583 21029
rect 5166 21020 5172 21032
rect 5224 21020 5230 21072
rect 5736 21060 5764 21100
rect 5902 21088 5908 21100
rect 5960 21088 5966 21140
rect 6914 21088 6920 21140
rect 6972 21128 6978 21140
rect 7561 21131 7619 21137
rect 7561 21128 7573 21131
rect 6972 21100 7573 21128
rect 6972 21088 6978 21100
rect 7561 21097 7573 21100
rect 7607 21097 7619 21131
rect 7561 21091 7619 21097
rect 8018 21088 8024 21140
rect 8076 21088 8082 21140
rect 8754 21088 8760 21140
rect 8812 21128 8818 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8812 21100 8953 21128
rect 8812 21088 8818 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 11882 21088 11888 21140
rect 11940 21088 11946 21140
rect 13078 21088 13084 21140
rect 13136 21088 13142 21140
rect 14366 21088 14372 21140
rect 14424 21088 14430 21140
rect 16393 21131 16451 21137
rect 16393 21097 16405 21131
rect 16439 21128 16451 21131
rect 17218 21128 17224 21140
rect 16439 21100 17224 21128
rect 16439 21097 16451 21100
rect 16393 21091 16451 21097
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 17865 21131 17923 21137
rect 17865 21097 17877 21131
rect 17911 21128 17923 21131
rect 17954 21128 17960 21140
rect 17911 21100 17960 21128
rect 17911 21097 17923 21100
rect 17865 21091 17923 21097
rect 17954 21088 17960 21100
rect 18012 21128 18018 21140
rect 18598 21128 18604 21140
rect 18012 21100 18604 21128
rect 18012 21088 18018 21100
rect 18598 21088 18604 21100
rect 18656 21088 18662 21140
rect 19702 21128 19708 21140
rect 19306 21100 19708 21128
rect 5460 21032 5764 21060
rect 1995 20964 2728 20992
rect 2777 20995 2835 21001
rect 1995 20961 2007 20964
rect 1949 20955 2007 20961
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 2866 20992 2872 21004
rect 2823 20964 2872 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 3326 20952 3332 21004
rect 3384 20992 3390 21004
rect 5460 20992 5488 21032
rect 7282 21020 7288 21072
rect 7340 21060 7346 21072
rect 7377 21063 7435 21069
rect 7377 21060 7389 21063
rect 7340 21032 7389 21060
rect 7340 21020 7346 21032
rect 7377 21029 7389 21032
rect 7423 21029 7435 21063
rect 7377 21023 7435 21029
rect 7466 21020 7472 21072
rect 7524 21060 7530 21072
rect 7524 21032 9536 21060
rect 7524 21020 7530 21032
rect 3384 20964 3556 20992
rect 3384 20952 3390 20964
rect 934 20884 940 20936
rect 992 20924 998 20936
rect 1397 20927 1455 20933
rect 1397 20924 1409 20927
rect 992 20896 1409 20924
rect 992 20884 998 20896
rect 1397 20893 1409 20896
rect 1443 20893 1455 20927
rect 1397 20887 1455 20893
rect 1857 20927 1915 20933
rect 1857 20893 1869 20927
rect 1903 20893 1915 20927
rect 1857 20887 1915 20893
rect 1872 20856 1900 20887
rect 2314 20884 2320 20936
rect 2372 20924 2378 20936
rect 2409 20927 2467 20933
rect 2409 20924 2421 20927
rect 2372 20896 2421 20924
rect 2372 20884 2378 20896
rect 2409 20893 2421 20896
rect 2455 20924 2467 20927
rect 3421 20927 3479 20933
rect 3421 20924 3433 20927
rect 2455 20896 3433 20924
rect 2455 20893 2467 20896
rect 2409 20887 2467 20893
rect 3421 20893 3433 20896
rect 3467 20893 3479 20927
rect 3528 20924 3556 20964
rect 4080 20964 5488 20992
rect 3970 20924 3976 20936
rect 3528 20896 3976 20924
rect 3421 20887 3479 20893
rect 3970 20884 3976 20896
rect 4028 20884 4034 20936
rect 4080 20933 4108 20964
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 5629 20995 5687 21001
rect 5629 20992 5641 20995
rect 5592 20964 5641 20992
rect 5592 20952 5598 20964
rect 5629 20961 5641 20964
rect 5675 20961 5687 20995
rect 5629 20955 5687 20961
rect 6638 20952 6644 21004
rect 6696 20992 6702 21004
rect 7745 20995 7803 21001
rect 7745 20992 7757 20995
rect 6696 20964 7757 20992
rect 6696 20952 6702 20964
rect 7745 20961 7757 20964
rect 7791 20961 7803 20995
rect 8205 20995 8263 21001
rect 8205 20992 8217 20995
rect 7745 20955 7803 20961
rect 7852 20964 8217 20992
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 4338 20884 4344 20936
rect 4396 20884 4402 20936
rect 4430 20884 4436 20936
rect 4488 20884 4494 20936
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20924 5227 20927
rect 5258 20924 5264 20936
rect 5215 20896 5264 20924
rect 5215 20893 5227 20896
rect 5169 20887 5227 20893
rect 5258 20884 5264 20896
rect 5316 20884 5322 20936
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20924 5411 20927
rect 7469 20927 7527 20933
rect 5399 20896 5672 20924
rect 5399 20893 5411 20896
rect 5353 20887 5411 20893
rect 3329 20859 3387 20865
rect 3329 20856 3341 20859
rect 1872 20828 3341 20856
rect 3329 20825 3341 20828
rect 3375 20825 3387 20859
rect 4448 20856 4476 20884
rect 4893 20859 4951 20865
rect 4893 20856 4905 20859
rect 4448 20828 4905 20856
rect 3329 20819 3387 20825
rect 4893 20825 4905 20828
rect 4939 20825 4951 20859
rect 5368 20856 5396 20887
rect 4893 20819 4951 20825
rect 5000 20828 5396 20856
rect 5644 20856 5672 20896
rect 7469 20893 7481 20927
rect 7515 20924 7527 20927
rect 7650 20924 7656 20936
rect 7515 20896 7656 20924
rect 7515 20893 7527 20896
rect 7469 20887 7527 20893
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 5810 20856 5816 20868
rect 5644 20828 5816 20856
rect 1578 20748 1584 20800
rect 1636 20748 1642 20800
rect 4249 20791 4307 20797
rect 4249 20757 4261 20791
rect 4295 20788 4307 20791
rect 5000 20788 5028 20828
rect 5810 20816 5816 20828
rect 5868 20816 5874 20868
rect 5902 20816 5908 20868
rect 5960 20816 5966 20868
rect 7852 20856 7880 20964
rect 8205 20961 8217 20964
rect 8251 20961 8263 20995
rect 8205 20955 8263 20961
rect 9398 20952 9404 21004
rect 9456 20952 9462 21004
rect 9508 21001 9536 21032
rect 14090 21020 14096 21072
rect 14148 21060 14154 21072
rect 19306 21060 19334 21100
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 21358 21088 21364 21140
rect 21416 21088 21422 21140
rect 14148 21032 19334 21060
rect 14148 21020 14154 21032
rect 9493 20995 9551 21001
rect 9493 20961 9505 20995
rect 9539 20961 9551 20995
rect 9493 20955 9551 20961
rect 11606 20952 11612 21004
rect 11664 20992 11670 21004
rect 15194 20992 15200 21004
rect 11664 20964 15200 20992
rect 11664 20952 11670 20964
rect 15194 20952 15200 20964
rect 15252 20992 15258 21004
rect 16114 20992 16120 21004
rect 15252 20964 16120 20992
rect 15252 20952 15258 20964
rect 16114 20952 16120 20964
rect 16172 20952 16178 21004
rect 16850 20992 16856 21004
rect 16224 20964 16856 20992
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 7130 20828 7880 20856
rect 4295 20760 5028 20788
rect 4295 20757 4307 20760
rect 4249 20751 4307 20757
rect 5534 20748 5540 20800
rect 5592 20748 5598 20800
rect 6730 20748 6736 20800
rect 6788 20788 6794 20800
rect 8128 20788 8156 20887
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 8720 20896 9321 20924
rect 8720 20884 8726 20896
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 12894 20884 12900 20936
rect 12952 20924 12958 20936
rect 12989 20927 13047 20933
rect 12989 20924 13001 20927
rect 12952 20896 13001 20924
rect 12952 20884 12958 20896
rect 12989 20893 13001 20896
rect 13035 20924 13047 20927
rect 13262 20924 13268 20936
rect 13035 20896 13268 20924
rect 13035 20893 13047 20896
rect 12989 20887 13047 20893
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 14274 20884 14280 20936
rect 14332 20884 14338 20936
rect 10413 20859 10471 20865
rect 10413 20825 10425 20859
rect 10459 20856 10471 20859
rect 10962 20856 10968 20868
rect 10459 20828 10968 20856
rect 10459 20825 10471 20828
rect 10413 20819 10471 20825
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 15838 20816 15844 20868
rect 15896 20856 15902 20868
rect 16224 20865 16252 20964
rect 16850 20952 16856 20964
rect 16908 20952 16914 21004
rect 19610 20952 19616 21004
rect 19668 20952 19674 21004
rect 22066 20964 23520 20992
rect 16574 20884 16580 20936
rect 16632 20884 16638 20936
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 17681 20927 17739 20933
rect 17681 20893 17693 20927
rect 17727 20924 17739 20927
rect 18046 20924 18052 20936
rect 17727 20896 18052 20924
rect 17727 20893 17739 20896
rect 17681 20887 17739 20893
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20924 21511 20927
rect 22066 20924 22094 20964
rect 23492 20936 23520 20964
rect 24026 20952 24032 21004
rect 24084 20992 24090 21004
rect 24084 20964 24532 20992
rect 24084 20952 24090 20964
rect 21499 20896 22094 20924
rect 23293 20927 23351 20933
rect 21499 20893 21511 20896
rect 21453 20887 21511 20893
rect 23293 20893 23305 20927
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 16209 20859 16267 20865
rect 16209 20856 16221 20859
rect 15896 20828 16221 20856
rect 15896 20816 15902 20828
rect 16209 20825 16221 20828
rect 16255 20825 16267 20859
rect 16209 20819 16267 20825
rect 16425 20859 16483 20865
rect 16425 20825 16437 20859
rect 16471 20856 16483 20859
rect 16592 20856 16620 20884
rect 17126 20856 17132 20868
rect 16471 20828 17132 20856
rect 16471 20825 16483 20828
rect 16425 20819 16483 20825
rect 17126 20816 17132 20828
rect 17184 20816 17190 20868
rect 19886 20816 19892 20868
rect 19944 20816 19950 20868
rect 21545 20859 21603 20865
rect 21545 20856 21557 20859
rect 21114 20828 21557 20856
rect 21545 20825 21557 20828
rect 21591 20825 21603 20859
rect 23308 20856 23336 20887
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 23845 20927 23903 20933
rect 23845 20924 23857 20927
rect 23532 20896 23857 20924
rect 23532 20884 23538 20896
rect 23845 20893 23857 20896
rect 23891 20924 23903 20927
rect 24302 20924 24308 20936
rect 23891 20896 24308 20924
rect 23891 20893 23903 20896
rect 23845 20887 23903 20893
rect 24302 20884 24308 20896
rect 24360 20884 24366 20936
rect 24504 20933 24532 20964
rect 24489 20927 24547 20933
rect 24489 20893 24501 20927
rect 24535 20924 24547 20927
rect 24762 20924 24768 20936
rect 24535 20896 24768 20924
rect 24535 20893 24547 20896
rect 24489 20887 24547 20893
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 25041 20859 25099 20865
rect 25041 20856 25053 20859
rect 23308 20828 25053 20856
rect 21545 20819 21603 20825
rect 25041 20825 25053 20828
rect 25087 20825 25099 20859
rect 25041 20819 25099 20825
rect 6788 20760 8156 20788
rect 6788 20748 6794 20760
rect 16574 20748 16580 20800
rect 16632 20748 16638 20800
rect 23382 20748 23388 20800
rect 23440 20748 23446 20800
rect 23937 20791 23995 20797
rect 23937 20757 23949 20791
rect 23983 20788 23995 20791
rect 24026 20788 24032 20800
rect 23983 20760 24032 20788
rect 23983 20757 23995 20760
rect 23937 20751 23995 20757
rect 24026 20748 24032 20760
rect 24084 20748 24090 20800
rect 1104 20698 26312 20720
rect 1104 20646 4761 20698
rect 4813 20646 4825 20698
rect 4877 20646 4889 20698
rect 4941 20646 4953 20698
rect 5005 20646 5017 20698
rect 5069 20646 11063 20698
rect 11115 20646 11127 20698
rect 11179 20646 11191 20698
rect 11243 20646 11255 20698
rect 11307 20646 11319 20698
rect 11371 20646 17365 20698
rect 17417 20646 17429 20698
rect 17481 20646 17493 20698
rect 17545 20646 17557 20698
rect 17609 20646 17621 20698
rect 17673 20646 23667 20698
rect 23719 20646 23731 20698
rect 23783 20646 23795 20698
rect 23847 20646 23859 20698
rect 23911 20646 23923 20698
rect 23975 20646 26312 20698
rect 1104 20624 26312 20646
rect 3418 20544 3424 20596
rect 3476 20544 3482 20596
rect 3973 20587 4031 20593
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 5258 20584 5264 20596
rect 4019 20556 5264 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 5258 20544 5264 20556
rect 5316 20584 5322 20596
rect 6914 20584 6920 20596
rect 5316 20556 6920 20584
rect 5316 20544 5322 20556
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 7466 20544 7472 20596
rect 7524 20544 7530 20596
rect 9306 20584 9312 20596
rect 8220 20556 9312 20584
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 2866 20448 2872 20460
rect 2823 20420 2872 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 2866 20408 2872 20420
rect 2924 20408 2930 20460
rect 3142 20408 3148 20460
rect 3200 20408 3206 20460
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 3436 20448 3464 20544
rect 5166 20476 5172 20528
rect 5224 20476 5230 20528
rect 5369 20519 5427 20525
rect 5369 20516 5381 20519
rect 5276 20488 5381 20516
rect 3605 20451 3663 20457
rect 3605 20448 3617 20451
rect 3283 20420 3372 20448
rect 3436 20420 3617 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 2884 20312 2912 20408
rect 3344 20312 3372 20420
rect 3605 20417 3617 20420
rect 3651 20417 3663 20451
rect 4338 20448 4344 20460
rect 3605 20411 3663 20417
rect 3712 20420 4344 20448
rect 3510 20340 3516 20392
rect 3568 20380 3574 20392
rect 3712 20389 3740 20420
rect 4338 20408 4344 20420
rect 4396 20448 4402 20460
rect 4617 20451 4675 20457
rect 4617 20448 4629 20451
rect 4396 20420 4629 20448
rect 4396 20408 4402 20420
rect 4617 20417 4629 20420
rect 4663 20417 4675 20451
rect 4617 20411 4675 20417
rect 4798 20408 4804 20460
rect 4856 20448 4862 20460
rect 5276 20448 5304 20488
rect 5369 20485 5381 20488
rect 5415 20485 5427 20519
rect 5369 20479 5427 20485
rect 6362 20476 6368 20528
rect 6420 20516 6426 20528
rect 8220 20516 8248 20556
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 10042 20544 10048 20596
rect 10100 20584 10106 20596
rect 10778 20584 10784 20596
rect 10100 20556 10784 20584
rect 10100 20544 10106 20556
rect 10778 20544 10784 20556
rect 10836 20584 10842 20596
rect 13173 20587 13231 20593
rect 13173 20584 13185 20587
rect 10836 20556 13185 20584
rect 10836 20544 10842 20556
rect 13173 20553 13185 20556
rect 13219 20553 13231 20587
rect 13173 20547 13231 20553
rect 19610 20544 19616 20596
rect 19668 20584 19674 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 19668 20556 19717 20584
rect 19668 20544 19674 20556
rect 19705 20553 19717 20556
rect 19751 20584 19763 20587
rect 19751 20556 22094 20584
rect 19751 20553 19763 20556
rect 19705 20547 19763 20553
rect 22066 20528 22094 20556
rect 6420 20488 8248 20516
rect 6420 20476 6426 20488
rect 4856 20420 5304 20448
rect 4856 20408 4862 20420
rect 5534 20408 5540 20460
rect 5592 20448 5598 20460
rect 5905 20451 5963 20457
rect 5905 20448 5917 20451
rect 5592 20420 5917 20448
rect 5592 20408 5598 20420
rect 5905 20417 5917 20420
rect 5951 20417 5963 20451
rect 5905 20411 5963 20417
rect 6270 20408 6276 20460
rect 6328 20448 6334 20460
rect 6546 20448 6552 20460
rect 6328 20420 6552 20448
rect 6328 20408 6334 20420
rect 6546 20408 6552 20420
rect 6604 20408 6610 20460
rect 8220 20457 8248 20488
rect 9214 20476 9220 20528
rect 9272 20476 9278 20528
rect 10134 20476 10140 20528
rect 10192 20516 10198 20528
rect 10597 20519 10655 20525
rect 10597 20516 10609 20519
rect 10192 20488 10609 20516
rect 10192 20476 10198 20488
rect 10597 20485 10609 20488
rect 10643 20485 10655 20519
rect 10597 20479 10655 20485
rect 10962 20476 10968 20528
rect 11020 20516 11026 20528
rect 12434 20516 12440 20528
rect 11020 20488 12440 20516
rect 11020 20476 11026 20488
rect 12434 20476 12440 20488
rect 12492 20476 12498 20528
rect 17037 20519 17095 20525
rect 17037 20485 17049 20519
rect 17083 20516 17095 20519
rect 17218 20516 17224 20528
rect 17083 20488 17224 20516
rect 17083 20485 17095 20488
rect 17037 20479 17095 20485
rect 17218 20476 17224 20488
rect 17276 20476 17282 20528
rect 17880 20488 20484 20516
rect 7101 20451 7159 20457
rect 7101 20448 7113 20451
rect 6656 20420 7113 20448
rect 3697 20383 3755 20389
rect 3697 20380 3709 20383
rect 3568 20352 3709 20380
rect 3568 20340 3574 20352
rect 3697 20349 3709 20352
rect 3743 20349 3755 20383
rect 3697 20343 3755 20349
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 5442 20380 5448 20392
rect 4755 20352 5448 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 5718 20340 5724 20392
rect 5776 20380 5782 20392
rect 6656 20380 6684 20420
rect 7101 20417 7113 20420
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 7285 20451 7343 20457
rect 7285 20417 7297 20451
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 11422 20448 11428 20460
rect 10551 20420 11428 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 5776 20352 6684 20380
rect 5776 20340 5782 20352
rect 6730 20340 6736 20392
rect 6788 20340 6794 20392
rect 6822 20340 6828 20392
rect 6880 20380 6886 20392
rect 7300 20380 7328 20411
rect 11422 20408 11428 20420
rect 11480 20408 11486 20460
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 6880 20352 7328 20380
rect 6880 20340 6886 20352
rect 8478 20340 8484 20392
rect 8536 20340 8542 20392
rect 10689 20383 10747 20389
rect 9508 20352 10548 20380
rect 5537 20315 5595 20321
rect 2884 20284 3280 20312
rect 3344 20284 4752 20312
rect 2866 20204 2872 20256
rect 2924 20204 2930 20256
rect 3252 20244 3280 20284
rect 4724 20256 4752 20284
rect 5537 20281 5549 20315
rect 5583 20312 5595 20315
rect 5583 20284 8340 20312
rect 5583 20281 5595 20284
rect 5537 20275 5595 20281
rect 3605 20247 3663 20253
rect 3605 20244 3617 20247
rect 3252 20216 3617 20244
rect 3605 20213 3617 20216
rect 3651 20244 3663 20247
rect 4430 20244 4436 20256
rect 3651 20216 4436 20244
rect 3651 20213 3663 20216
rect 3605 20207 3663 20213
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 4522 20204 4528 20256
rect 4580 20244 4586 20256
rect 4617 20247 4675 20253
rect 4617 20244 4629 20247
rect 4580 20216 4629 20244
rect 4580 20204 4586 20216
rect 4617 20213 4629 20216
rect 4663 20213 4675 20247
rect 4617 20207 4675 20213
rect 4706 20204 4712 20256
rect 4764 20244 4770 20256
rect 4985 20247 5043 20253
rect 4985 20244 4997 20247
rect 4764 20216 4997 20244
rect 4764 20204 4770 20216
rect 4985 20213 4997 20216
rect 5031 20213 5043 20247
rect 4985 20207 5043 20213
rect 5350 20204 5356 20256
rect 5408 20204 5414 20256
rect 6086 20204 6092 20256
rect 6144 20204 6150 20256
rect 6270 20204 6276 20256
rect 6328 20244 6334 20256
rect 6730 20244 6736 20256
rect 6328 20216 6736 20244
rect 6328 20204 6334 20216
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 8312 20244 8340 20284
rect 9508 20244 9536 20352
rect 9582 20272 9588 20324
rect 9640 20312 9646 20324
rect 10137 20315 10195 20321
rect 10137 20312 10149 20315
rect 9640 20284 10149 20312
rect 9640 20272 9646 20284
rect 10137 20281 10149 20284
rect 10183 20281 10195 20315
rect 10520 20312 10548 20352
rect 10689 20349 10701 20383
rect 10735 20349 10747 20383
rect 13004 20380 13032 20411
rect 13446 20408 13452 20460
rect 13504 20408 13510 20460
rect 13630 20408 13636 20460
rect 13688 20408 13694 20460
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 15252 20420 15761 20448
rect 15252 20408 15258 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 16850 20408 16856 20460
rect 16908 20408 16914 20460
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 17880 20457 17908 20488
rect 20456 20460 20484 20488
rect 22002 20476 22008 20528
rect 22060 20516 22094 20528
rect 22060 20488 22968 20516
rect 22060 20476 22066 20488
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 17954 20408 17960 20460
rect 18012 20408 18018 20460
rect 18233 20451 18291 20457
rect 18233 20417 18245 20451
rect 18279 20448 18291 20451
rect 19058 20448 19064 20460
rect 18279 20420 19064 20448
rect 18279 20417 18291 20420
rect 18233 20411 18291 20417
rect 19058 20408 19064 20420
rect 19116 20408 19122 20460
rect 20438 20408 20444 20460
rect 20496 20448 20502 20460
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 20496 20420 20545 20448
rect 20496 20408 20502 20420
rect 20533 20417 20545 20420
rect 20579 20448 20591 20451
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20579 20420 21005 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20993 20417 21005 20420
rect 21039 20448 21051 20451
rect 21450 20448 21456 20460
rect 21039 20420 21456 20448
rect 21039 20417 21051 20420
rect 20993 20411 21051 20417
rect 21450 20408 21456 20420
rect 21508 20408 21514 20460
rect 22940 20457 22968 20488
rect 24026 20476 24032 20528
rect 24084 20476 24090 20528
rect 24762 20476 24768 20528
rect 24820 20476 24826 20528
rect 22925 20451 22983 20457
rect 22925 20417 22937 20451
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20448 23351 20451
rect 23382 20448 23388 20460
rect 23339 20420 23388 20448
rect 23339 20417 23351 20420
rect 23293 20411 23351 20417
rect 23382 20408 23388 20420
rect 23440 20408 23446 20460
rect 13817 20383 13875 20389
rect 13817 20380 13829 20383
rect 13004 20352 13829 20380
rect 10689 20343 10747 20349
rect 13817 20349 13829 20352
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 13924 20352 16160 20380
rect 10704 20312 10732 20343
rect 10520 20284 10732 20312
rect 10137 20275 10195 20281
rect 13262 20272 13268 20324
rect 13320 20312 13326 20324
rect 13924 20312 13952 20352
rect 13320 20284 13952 20312
rect 15565 20315 15623 20321
rect 13320 20272 13326 20284
rect 15565 20281 15577 20315
rect 15611 20312 15623 20315
rect 16132 20312 16160 20352
rect 17770 20340 17776 20392
rect 17828 20380 17834 20392
rect 18141 20383 18199 20389
rect 18141 20380 18153 20383
rect 17828 20352 18153 20380
rect 17828 20340 17834 20352
rect 18141 20349 18153 20352
rect 18187 20349 18199 20383
rect 18141 20343 18199 20349
rect 20622 20340 20628 20392
rect 20680 20340 20686 20392
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 20956 20352 21281 20380
rect 20956 20340 20962 20352
rect 21269 20349 21281 20352
rect 21315 20380 21327 20383
rect 21634 20380 21640 20392
rect 21315 20352 21640 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 25130 20380 25136 20392
rect 22066 20352 25136 20380
rect 15611 20284 16068 20312
rect 16132 20284 18184 20312
rect 15611 20281 15623 20284
rect 15565 20275 15623 20281
rect 16040 20256 16068 20284
rect 8312 20216 9536 20244
rect 9950 20204 9956 20256
rect 10008 20204 10014 20256
rect 15657 20247 15715 20253
rect 15657 20213 15669 20247
rect 15703 20244 15715 20247
rect 15930 20244 15936 20256
rect 15703 20216 15936 20244
rect 15703 20213 15715 20216
rect 15657 20207 15715 20213
rect 15930 20204 15936 20216
rect 15988 20204 15994 20256
rect 16022 20204 16028 20256
rect 16080 20204 16086 20256
rect 16209 20247 16267 20253
rect 16209 20213 16221 20247
rect 16255 20244 16267 20247
rect 16298 20244 16304 20256
rect 16255 20216 16304 20244
rect 16255 20213 16267 20216
rect 16209 20207 16267 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16632 20216 16681 20244
rect 16632 20204 16638 20216
rect 16669 20213 16681 20216
rect 16715 20213 16727 20247
rect 16669 20207 16727 20213
rect 18046 20204 18052 20256
rect 18104 20204 18110 20256
rect 18156 20244 18184 20284
rect 18230 20272 18236 20324
rect 18288 20312 18294 20324
rect 22066 20312 22094 20352
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 18288 20284 22094 20312
rect 18288 20272 18294 20284
rect 18506 20244 18512 20256
rect 18156 20216 18512 20244
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 20809 20247 20867 20253
rect 20809 20213 20821 20247
rect 20855 20244 20867 20247
rect 20990 20244 20996 20256
rect 20855 20216 20996 20244
rect 20855 20213 20867 20216
rect 20809 20207 20867 20213
rect 20990 20204 20996 20216
rect 21048 20204 21054 20256
rect 21266 20204 21272 20256
rect 21324 20204 21330 20256
rect 21358 20204 21364 20256
rect 21416 20244 21422 20256
rect 21545 20247 21603 20253
rect 21545 20244 21557 20247
rect 21416 20216 21557 20244
rect 21416 20204 21422 20216
rect 21545 20213 21557 20216
rect 21591 20213 21603 20247
rect 21545 20207 21603 20213
rect 1104 20154 26312 20176
rect 1104 20102 4101 20154
rect 4153 20102 4165 20154
rect 4217 20102 4229 20154
rect 4281 20102 4293 20154
rect 4345 20102 4357 20154
rect 4409 20102 10403 20154
rect 10455 20102 10467 20154
rect 10519 20102 10531 20154
rect 10583 20102 10595 20154
rect 10647 20102 10659 20154
rect 10711 20102 16705 20154
rect 16757 20102 16769 20154
rect 16821 20102 16833 20154
rect 16885 20102 16897 20154
rect 16949 20102 16961 20154
rect 17013 20102 23007 20154
rect 23059 20102 23071 20154
rect 23123 20102 23135 20154
rect 23187 20102 23199 20154
rect 23251 20102 23263 20154
rect 23315 20102 26312 20154
rect 1104 20080 26312 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2924 20012 2973 20040
rect 2924 20000 2930 20012
rect 2961 20009 2973 20012
rect 3007 20040 3019 20043
rect 3418 20040 3424 20052
rect 3007 20012 3424 20040
rect 3007 20009 3019 20012
rect 2961 20003 3019 20009
rect 3418 20000 3424 20012
rect 3476 20000 3482 20052
rect 4430 20000 4436 20052
rect 4488 20000 4494 20052
rect 4617 20043 4675 20049
rect 4617 20009 4629 20043
rect 4663 20040 4675 20043
rect 4798 20040 4804 20052
rect 4663 20012 4804 20040
rect 4663 20009 4675 20012
rect 4617 20003 4675 20009
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 4985 20043 5043 20049
rect 4985 20009 4997 20043
rect 5031 20040 5043 20043
rect 5350 20040 5356 20052
rect 5031 20012 5356 20040
rect 5031 20009 5043 20012
rect 4985 20003 5043 20009
rect 4448 19972 4476 20000
rect 5000 19972 5028 20003
rect 5350 20000 5356 20012
rect 5408 20000 5414 20052
rect 5718 20000 5724 20052
rect 5776 20000 5782 20052
rect 5902 20000 5908 20052
rect 5960 20000 5966 20052
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7009 20043 7067 20049
rect 7009 20040 7021 20043
rect 6972 20012 7021 20040
rect 6972 20000 6978 20012
rect 7009 20009 7021 20012
rect 7055 20009 7067 20043
rect 7009 20003 7067 20009
rect 9214 20000 9220 20052
rect 9272 20000 9278 20052
rect 9950 20040 9956 20052
rect 9784 20012 9956 20040
rect 4448 19944 5028 19972
rect 6362 19932 6368 19984
rect 6420 19972 6426 19984
rect 6638 19972 6644 19984
rect 6420 19944 6644 19972
rect 6420 19932 6426 19944
rect 6638 19932 6644 19944
rect 6696 19972 6702 19984
rect 6733 19975 6791 19981
rect 6733 19972 6745 19975
rect 6696 19944 6745 19972
rect 6696 19932 6702 19944
rect 6733 19941 6745 19944
rect 6779 19941 6791 19975
rect 6733 19935 6791 19941
rect 7469 19975 7527 19981
rect 7469 19941 7481 19975
rect 7515 19972 7527 19975
rect 9784 19972 9812 20012
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 11422 20000 11428 20052
rect 11480 20000 11486 20052
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 12342 20040 12348 20052
rect 11756 20012 12348 20040
rect 11756 20000 11762 20012
rect 12342 20000 12348 20012
rect 12400 20040 12406 20052
rect 12713 20043 12771 20049
rect 12713 20040 12725 20043
rect 12400 20012 12725 20040
rect 12400 20000 12406 20012
rect 12713 20009 12725 20012
rect 12759 20009 12771 20043
rect 12713 20003 12771 20009
rect 15948 20012 16804 20040
rect 7515 19944 8616 19972
rect 7515 19941 7527 19944
rect 7469 19935 7527 19941
rect 3510 19904 3516 19916
rect 2424 19876 2728 19904
rect 2424 19845 2452 19876
rect 2409 19839 2467 19845
rect 2409 19805 2421 19839
rect 2455 19805 2467 19839
rect 2409 19799 2467 19805
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19805 2651 19839
rect 2593 19799 2651 19805
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2501 19703 2559 19709
rect 2501 19700 2513 19703
rect 1728 19672 2513 19700
rect 1728 19660 1734 19672
rect 2501 19669 2513 19672
rect 2547 19669 2559 19703
rect 2608 19700 2636 19799
rect 2700 19768 2728 19876
rect 2976 19876 3516 19904
rect 2976 19848 3004 19876
rect 3510 19864 3516 19876
rect 3568 19864 3574 19916
rect 3605 19907 3663 19913
rect 3605 19873 3617 19907
rect 3651 19904 3663 19907
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3651 19876 4445 19904
rect 3651 19873 3663 19876
rect 3605 19867 3663 19873
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 5166 19864 5172 19916
rect 5224 19864 5230 19916
rect 5442 19864 5448 19916
rect 5500 19904 5506 19916
rect 7098 19904 7104 19916
rect 5500 19876 7104 19904
rect 5500 19864 5506 19876
rect 2774 19796 2780 19848
rect 2832 19796 2838 19848
rect 2958 19796 2964 19848
rect 3016 19796 3022 19848
rect 3326 19796 3332 19848
rect 3384 19796 3390 19848
rect 3418 19796 3424 19848
rect 3476 19796 3482 19848
rect 3528 19836 3556 19864
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 3528 19808 3801 19836
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19836 4583 19839
rect 4706 19836 4712 19848
rect 4571 19808 4712 19836
rect 4571 19805 4583 19808
rect 4525 19799 4583 19805
rect 3605 19771 3663 19777
rect 3605 19768 3617 19771
rect 2700 19740 3617 19768
rect 3605 19737 3617 19740
rect 3651 19737 3663 19771
rect 3804 19768 3832 19799
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19805 4951 19839
rect 4893 19799 4951 19805
rect 5629 19839 5687 19845
rect 5629 19805 5641 19839
rect 5675 19836 5687 19839
rect 5718 19836 5724 19848
rect 5675 19808 5724 19836
rect 5675 19805 5687 19808
rect 5629 19799 5687 19805
rect 4908 19768 4936 19799
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5810 19796 5816 19848
rect 5868 19796 5874 19848
rect 6086 19796 6092 19848
rect 6144 19796 6150 19848
rect 6196 19845 6224 19876
rect 6932 19845 6960 19876
rect 7098 19864 7104 19876
rect 7156 19904 7162 19916
rect 7650 19904 7656 19916
rect 7156 19876 7656 19904
rect 7156 19864 7162 19876
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 8588 19913 8616 19944
rect 9048 19944 9812 19972
rect 11440 19972 11468 20000
rect 12618 19972 12624 19984
rect 11440 19944 12624 19972
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 6564 19768 6592 19799
rect 7282 19796 7288 19848
rect 7340 19796 7346 19848
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19836 8539 19839
rect 9048 19836 9076 19944
rect 12618 19932 12624 19944
rect 12676 19932 12682 19984
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9364 19876 9689 19904
rect 9364 19864 9370 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 13630 19864 13636 19916
rect 13688 19904 13694 19916
rect 13688 19876 14320 19904
rect 13688 19864 13694 19876
rect 8527 19808 9076 19836
rect 8527 19805 8539 19808
rect 8481 19799 8539 19805
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9582 19796 9588 19848
rect 9640 19796 9646 19848
rect 11422 19836 11428 19848
rect 11086 19808 11428 19836
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19805 12587 19839
rect 12529 19799 12587 19805
rect 6638 19768 6644 19780
rect 3804 19740 4936 19768
rect 5000 19740 6644 19768
rect 3605 19731 3663 19737
rect 3145 19703 3203 19709
rect 3145 19700 3157 19703
rect 2608 19672 3157 19700
rect 2501 19663 2559 19669
rect 3145 19669 3157 19672
rect 3191 19700 3203 19703
rect 4430 19700 4436 19712
rect 3191 19672 4436 19700
rect 3191 19669 3203 19672
rect 3145 19663 3203 19669
rect 4430 19660 4436 19672
rect 4488 19660 4494 19712
rect 4522 19660 4528 19712
rect 4580 19700 4586 19712
rect 5000 19700 5028 19740
rect 6638 19728 6644 19740
rect 6696 19768 6702 19780
rect 7300 19768 7328 19796
rect 6696 19740 7328 19768
rect 6696 19728 6702 19740
rect 7926 19728 7932 19780
rect 7984 19768 7990 19780
rect 8389 19771 8447 19777
rect 8389 19768 8401 19771
rect 7984 19740 8401 19768
rect 7984 19728 7990 19740
rect 8389 19737 8401 19740
rect 8435 19737 8447 19771
rect 9953 19771 10011 19777
rect 9953 19768 9965 19771
rect 8389 19731 8447 19737
rect 9416 19740 9965 19768
rect 4580 19672 5028 19700
rect 4580 19660 4586 19672
rect 5350 19660 5356 19712
rect 5408 19700 5414 19712
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 5408 19672 5457 19700
rect 5408 19660 5414 19672
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 5445 19663 5503 19669
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 6365 19703 6423 19709
rect 6365 19700 6377 19703
rect 6052 19672 6377 19700
rect 6052 19660 6058 19672
rect 6365 19669 6377 19672
rect 6411 19700 6423 19703
rect 6730 19700 6736 19712
rect 6411 19672 6736 19700
rect 6411 19669 6423 19672
rect 6365 19663 6423 19669
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 8018 19660 8024 19712
rect 8076 19660 8082 19712
rect 9416 19709 9444 19740
rect 9953 19737 9965 19740
rect 9999 19737 10011 19771
rect 12544 19768 12572 19799
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 12805 19839 12863 19845
rect 12805 19836 12817 19839
rect 12768 19808 12817 19836
rect 12768 19796 12774 19808
rect 12805 19805 12817 19808
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 14292 19845 14320 19876
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 13504 19808 14105 19836
rect 13504 19796 13510 19808
rect 14093 19805 14105 19808
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 13998 19768 14004 19780
rect 12544 19740 14004 19768
rect 9953 19731 10011 19737
rect 13998 19728 14004 19740
rect 14056 19728 14062 19780
rect 14108 19768 14136 19799
rect 15948 19768 15976 20012
rect 16482 19972 16488 19984
rect 16040 19944 16488 19972
rect 16040 19845 16068 19944
rect 16482 19932 16488 19944
rect 16540 19932 16546 19984
rect 16574 19932 16580 19984
rect 16632 19972 16638 19984
rect 16776 19972 16804 20012
rect 19886 20000 19892 20052
rect 19944 20040 19950 20052
rect 20073 20043 20131 20049
rect 20073 20040 20085 20043
rect 19944 20012 20085 20040
rect 19944 20000 19950 20012
rect 20073 20009 20085 20012
rect 20119 20009 20131 20043
rect 25958 20040 25964 20052
rect 20073 20003 20131 20009
rect 20180 20012 25964 20040
rect 20180 19972 20208 20012
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 21818 19972 21824 19984
rect 16632 19944 16712 19972
rect 16776 19944 20208 19972
rect 20272 19944 21824 19972
rect 16632 19932 16638 19944
rect 16316 19876 16620 19904
rect 16316 19848 16344 19876
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19805 16083 19839
rect 16025 19799 16083 19805
rect 16298 19796 16304 19848
rect 16356 19796 16362 19848
rect 16482 19796 16488 19848
rect 16540 19796 16546 19848
rect 16592 19845 16620 19876
rect 16684 19845 16712 19944
rect 19426 19864 19432 19916
rect 19484 19864 19490 19916
rect 16577 19839 16635 19845
rect 16577 19805 16589 19839
rect 16623 19805 16635 19839
rect 16577 19799 16635 19805
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 14108 19740 15976 19768
rect 16209 19771 16267 19777
rect 16209 19737 16221 19771
rect 16255 19768 16267 19771
rect 16684 19768 16712 19799
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19836 18107 19839
rect 18230 19836 18236 19848
rect 18095 19808 18236 19836
rect 18095 19805 18107 19808
rect 18049 19799 18107 19805
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19208 19808 19257 19836
rect 19208 19796 19214 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 20162 19796 20168 19848
rect 20220 19836 20226 19848
rect 20272 19845 20300 19944
rect 21818 19932 21824 19944
rect 21876 19932 21882 19984
rect 20438 19864 20444 19916
rect 20496 19864 20502 19916
rect 20990 19864 20996 19916
rect 21048 19904 21054 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 21048 19876 21741 19904
rect 21048 19864 21054 19876
rect 21729 19873 21741 19876
rect 21775 19873 21787 19907
rect 21729 19867 21787 19873
rect 22002 19864 22008 19916
rect 22060 19864 22066 19916
rect 22278 19864 22284 19916
rect 22336 19904 22342 19916
rect 24029 19907 24087 19913
rect 24029 19904 24041 19907
rect 22336 19876 24041 19904
rect 22336 19864 22342 19876
rect 24029 19873 24041 19876
rect 24075 19873 24087 19907
rect 24029 19867 24087 19873
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 20220 19808 20269 19836
rect 20220 19796 20226 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 20395 19808 20484 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 20456 19780 20484 19808
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 20809 19839 20867 19845
rect 20809 19805 20821 19839
rect 20855 19805 20867 19839
rect 20809 19799 20867 19805
rect 16255 19740 16712 19768
rect 16255 19737 16267 19740
rect 16209 19731 16267 19737
rect 20438 19728 20444 19780
rect 20496 19768 20502 19780
rect 20824 19768 20852 19799
rect 21266 19796 21272 19848
rect 21324 19796 21330 19848
rect 21358 19796 21364 19848
rect 21416 19796 21422 19848
rect 20496 19740 20852 19768
rect 20496 19728 20502 19740
rect 21174 19728 21180 19780
rect 21232 19768 21238 19780
rect 21453 19771 21511 19777
rect 21453 19768 21465 19771
rect 21232 19740 21465 19768
rect 21232 19728 21238 19740
rect 21453 19737 21465 19740
rect 21499 19737 21511 19771
rect 21453 19731 21511 19737
rect 21542 19728 21548 19780
rect 21600 19777 21606 19780
rect 21600 19771 21629 19777
rect 21617 19737 21629 19771
rect 21600 19731 21629 19737
rect 22281 19771 22339 19777
rect 22281 19737 22293 19771
rect 22327 19737 22339 19771
rect 22281 19731 22339 19737
rect 21600 19728 21606 19731
rect 9401 19703 9459 19709
rect 9401 19669 9413 19703
rect 9447 19669 9459 19703
rect 9401 19663 9459 19669
rect 12802 19660 12808 19712
rect 12860 19700 12866 19712
rect 12897 19703 12955 19709
rect 12897 19700 12909 19703
rect 12860 19672 12909 19700
rect 12860 19660 12866 19672
rect 12897 19669 12909 19672
rect 12943 19669 12955 19703
rect 12897 19663 12955 19669
rect 14090 19660 14096 19712
rect 14148 19700 14154 19712
rect 14185 19703 14243 19709
rect 14185 19700 14197 19703
rect 14148 19672 14197 19700
rect 14148 19660 14154 19672
rect 14185 19669 14197 19672
rect 14231 19669 14243 19703
rect 14185 19663 14243 19669
rect 15841 19703 15899 19709
rect 15841 19669 15853 19703
rect 15887 19700 15899 19703
rect 16114 19700 16120 19712
rect 15887 19672 16120 19700
rect 15887 19669 15899 19672
rect 15841 19663 15899 19669
rect 16114 19660 16120 19672
rect 16172 19660 16178 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 16853 19703 16911 19709
rect 16853 19700 16865 19703
rect 16632 19672 16865 19700
rect 16632 19660 16638 19672
rect 16853 19669 16865 19672
rect 16899 19669 16911 19703
rect 16853 19663 16911 19669
rect 17770 19660 17776 19712
rect 17828 19700 17834 19712
rect 18233 19703 18291 19709
rect 18233 19700 18245 19703
rect 17828 19672 18245 19700
rect 17828 19660 17834 19672
rect 18233 19669 18245 19672
rect 18279 19669 18291 19703
rect 18233 19663 18291 19669
rect 20898 19660 20904 19712
rect 20956 19660 20962 19712
rect 21085 19703 21143 19709
rect 21085 19669 21097 19703
rect 21131 19700 21143 19703
rect 22296 19700 22324 19731
rect 23290 19728 23296 19780
rect 23348 19728 23354 19780
rect 21131 19672 22324 19700
rect 21131 19669 21143 19672
rect 21085 19663 21143 19669
rect 1104 19610 26312 19632
rect 1104 19558 4761 19610
rect 4813 19558 4825 19610
rect 4877 19558 4889 19610
rect 4941 19558 4953 19610
rect 5005 19558 5017 19610
rect 5069 19558 11063 19610
rect 11115 19558 11127 19610
rect 11179 19558 11191 19610
rect 11243 19558 11255 19610
rect 11307 19558 11319 19610
rect 11371 19558 17365 19610
rect 17417 19558 17429 19610
rect 17481 19558 17493 19610
rect 17545 19558 17557 19610
rect 17609 19558 17621 19610
rect 17673 19558 23667 19610
rect 23719 19558 23731 19610
rect 23783 19558 23795 19610
rect 23847 19558 23859 19610
rect 23911 19558 23923 19610
rect 23975 19558 26312 19610
rect 1104 19536 26312 19558
rect 2958 19456 2964 19508
rect 3016 19496 3022 19508
rect 3145 19499 3203 19505
rect 3145 19496 3157 19499
rect 3016 19468 3157 19496
rect 3016 19456 3022 19468
rect 3145 19465 3157 19468
rect 3191 19465 3203 19499
rect 3145 19459 3203 19465
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 4488 19468 4752 19496
rect 4488 19456 4494 19468
rect 1670 19388 1676 19440
rect 1728 19388 1734 19440
rect 4614 19428 4620 19440
rect 3804 19400 4620 19428
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 3804 19369 3832 19400
rect 4614 19388 4620 19400
rect 4672 19388 4678 19440
rect 4724 19428 4752 19468
rect 4798 19456 4804 19508
rect 4856 19456 4862 19508
rect 8389 19499 8447 19505
rect 8389 19465 8401 19499
rect 8435 19496 8447 19499
rect 8478 19496 8484 19508
rect 8435 19468 8484 19496
rect 8435 19465 8447 19468
rect 8389 19459 8447 19465
rect 8478 19456 8484 19468
rect 8536 19456 8542 19508
rect 12710 19496 12716 19508
rect 11716 19468 12716 19496
rect 7190 19428 7196 19440
rect 4724 19400 7196 19428
rect 7190 19388 7196 19400
rect 7248 19388 7254 19440
rect 9306 19388 9312 19440
rect 9364 19428 9370 19440
rect 11609 19431 11667 19437
rect 11609 19428 11621 19431
rect 9364 19400 9628 19428
rect 11086 19400 11621 19428
rect 9364 19388 9370 19400
rect 3237 19363 3295 19369
rect 3237 19329 3249 19363
rect 3283 19360 3295 19363
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 3283 19332 3801 19360
rect 3283 19329 3295 19332
rect 3237 19323 3295 19329
rect 3789 19329 3801 19332
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19360 4031 19363
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 4019 19332 4261 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4249 19329 4261 19332
rect 4295 19360 4307 19363
rect 5166 19360 5172 19372
rect 4295 19332 5172 19360
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3329 19295 3387 19301
rect 3329 19292 3341 19295
rect 3200 19264 3341 19292
rect 3200 19252 3206 19264
rect 3329 19261 3341 19264
rect 3375 19292 3387 19295
rect 3988 19292 4016 19323
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 5810 19320 5816 19372
rect 5868 19360 5874 19372
rect 6362 19360 6368 19372
rect 5868 19332 6368 19360
rect 5868 19320 5874 19332
rect 6362 19320 6368 19332
rect 6420 19320 6426 19372
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 6730 19360 6736 19372
rect 6595 19332 6736 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 6730 19320 6736 19332
rect 6788 19320 6794 19372
rect 8018 19320 8024 19372
rect 8076 19360 8082 19372
rect 8573 19363 8631 19369
rect 8573 19360 8585 19363
rect 8076 19332 8585 19360
rect 8076 19320 8082 19332
rect 8573 19329 8585 19332
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 9600 19369 9628 19400
rect 11609 19397 11621 19400
rect 11655 19397 11667 19431
rect 11609 19391 11667 19397
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 11716 19360 11744 19468
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 13541 19499 13599 19505
rect 13541 19465 13553 19499
rect 13587 19496 13599 19499
rect 13833 19499 13891 19505
rect 13833 19496 13845 19499
rect 13587 19468 13845 19496
rect 13587 19465 13599 19468
rect 13541 19459 13599 19465
rect 13833 19465 13845 19468
rect 13879 19465 13891 19499
rect 13833 19459 13891 19465
rect 13998 19456 14004 19508
rect 14056 19456 14062 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 16393 19499 16451 19505
rect 16393 19496 16405 19499
rect 15252 19468 16405 19496
rect 15252 19456 15258 19468
rect 16393 19465 16405 19468
rect 16439 19465 16451 19499
rect 16393 19459 16451 19465
rect 17037 19499 17095 19505
rect 17037 19465 17049 19499
rect 17083 19496 17095 19499
rect 18141 19499 18199 19505
rect 18141 19496 18153 19499
rect 17083 19468 18153 19496
rect 17083 19465 17095 19468
rect 17037 19459 17095 19465
rect 18141 19465 18153 19468
rect 18187 19465 18199 19499
rect 18141 19459 18199 19465
rect 20257 19499 20315 19505
rect 20257 19465 20269 19499
rect 20303 19465 20315 19499
rect 20257 19459 20315 19465
rect 20349 19499 20407 19505
rect 20349 19465 20361 19499
rect 20395 19496 20407 19499
rect 20530 19496 20536 19508
rect 20395 19468 20536 19496
rect 20395 19465 20407 19468
rect 20349 19459 20407 19465
rect 12066 19428 12072 19440
rect 11808 19400 12072 19428
rect 11808 19369 11836 19400
rect 12066 19388 12072 19400
rect 12124 19388 12130 19440
rect 12802 19388 12808 19440
rect 12860 19388 12866 19440
rect 13630 19388 13636 19440
rect 13688 19388 13694 19440
rect 17512 19400 17724 19428
rect 11572 19332 11744 19360
rect 11793 19363 11851 19369
rect 11572 19320 11578 19332
rect 11793 19329 11805 19363
rect 11839 19329 11851 19363
rect 11793 19323 11851 19329
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19329 15899 19363
rect 15841 19323 15899 19329
rect 4338 19292 4344 19304
rect 3375 19264 4016 19292
rect 4080 19264 4344 19292
rect 3375 19261 3387 19264
rect 3329 19255 3387 19261
rect 3418 19116 3424 19168
rect 3476 19116 3482 19168
rect 3602 19116 3608 19168
rect 3660 19116 3666 19168
rect 3973 19159 4031 19165
rect 3973 19125 3985 19159
rect 4019 19156 4031 19159
rect 4080 19156 4108 19264
rect 4338 19252 4344 19264
rect 4396 19292 4402 19304
rect 4525 19295 4583 19301
rect 4525 19292 4537 19295
rect 4396 19264 4537 19292
rect 4396 19252 4402 19264
rect 4525 19261 4537 19264
rect 4571 19261 4583 19295
rect 9861 19295 9919 19301
rect 9861 19292 9873 19295
rect 4525 19255 4583 19261
rect 9692 19264 9873 19292
rect 4157 19227 4215 19233
rect 4157 19193 4169 19227
rect 4203 19224 4215 19227
rect 4430 19224 4436 19236
rect 4203 19196 4436 19224
rect 4203 19193 4215 19196
rect 4157 19187 4215 19193
rect 4430 19184 4436 19196
rect 4488 19184 4494 19236
rect 9309 19227 9367 19233
rect 9309 19193 9321 19227
rect 9355 19224 9367 19227
rect 9692 19224 9720 19264
rect 9861 19261 9873 19264
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 12069 19295 12127 19301
rect 12069 19261 12081 19295
rect 12115 19292 12127 19295
rect 12158 19292 12164 19304
rect 12115 19264 12164 19292
rect 12115 19261 12127 19264
rect 12069 19255 12127 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 15746 19252 15752 19304
rect 15804 19252 15810 19304
rect 15856 19292 15884 19323
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 15988 19332 16221 19360
rect 15988 19320 15994 19332
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17512 19369 17540 19400
rect 17497 19363 17555 19369
rect 17184 19332 17448 19360
rect 17184 19320 17190 19332
rect 17218 19292 17224 19304
rect 15856 19264 17224 19292
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17420 19292 17448 19332
rect 17497 19329 17509 19363
rect 17543 19329 17555 19363
rect 17497 19323 17555 19329
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19329 17647 19363
rect 17696 19360 17724 19400
rect 17862 19388 17868 19440
rect 17920 19388 17926 19440
rect 17954 19388 17960 19440
rect 18012 19428 18018 19440
rect 18877 19431 18935 19437
rect 18877 19428 18889 19431
rect 18012 19400 18889 19428
rect 18012 19388 18018 19400
rect 18877 19397 18889 19400
rect 18923 19397 18935 19431
rect 19150 19428 19156 19440
rect 18877 19391 18935 19397
rect 18984 19400 19156 19428
rect 18046 19360 18052 19372
rect 17696 19332 18052 19360
rect 17589 19323 17647 19329
rect 17604 19292 17632 19323
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 18138 19320 18144 19372
rect 18196 19360 18202 19372
rect 18233 19363 18291 19369
rect 18233 19360 18245 19363
rect 18196 19332 18245 19360
rect 18196 19320 18202 19332
rect 18233 19329 18245 19332
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18984 19360 19012 19400
rect 19150 19388 19156 19400
rect 19208 19388 19214 19440
rect 19889 19431 19947 19437
rect 19889 19397 19901 19431
rect 19935 19428 19947 19431
rect 19978 19428 19984 19440
rect 19935 19400 19984 19428
rect 19935 19397 19947 19400
rect 19889 19391 19947 19397
rect 19978 19388 19984 19400
rect 20036 19388 20042 19440
rect 20162 19437 20168 19440
rect 20105 19431 20168 19437
rect 20105 19397 20117 19431
rect 20151 19397 20168 19431
rect 20105 19391 20168 19397
rect 20162 19388 20168 19391
rect 20220 19388 20226 19440
rect 20272 19428 20300 19459
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 21266 19456 21272 19508
rect 21324 19496 21330 19508
rect 22189 19499 22247 19505
rect 22189 19496 22201 19499
rect 21324 19468 22201 19496
rect 21324 19456 21330 19468
rect 22189 19465 22201 19468
rect 22235 19465 22247 19499
rect 22189 19459 22247 19465
rect 23201 19499 23259 19505
rect 23201 19465 23213 19499
rect 23247 19496 23259 19499
rect 23290 19496 23296 19508
rect 23247 19468 23296 19496
rect 23247 19465 23259 19468
rect 23201 19459 23259 19465
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 20714 19428 20720 19440
rect 20272 19400 20720 19428
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 20898 19388 20904 19440
rect 20956 19428 20962 19440
rect 20956 19400 21496 19428
rect 20956 19388 20962 19400
rect 18371 19332 19012 19360
rect 19061 19363 19119 19369
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 19061 19329 19073 19363
rect 19107 19360 19119 19363
rect 19334 19360 19340 19372
rect 19107 19332 19340 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 20523 19363 20581 19369
rect 20523 19329 20535 19363
rect 20569 19329 20581 19363
rect 20523 19323 20581 19329
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 21082 19360 21088 19372
rect 20855 19332 21088 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 17420 19264 17632 19292
rect 16574 19224 16580 19236
rect 9355 19196 9720 19224
rect 16224 19196 16580 19224
rect 9355 19193 9367 19196
rect 9309 19187 9367 19193
rect 4019 19128 4108 19156
rect 4019 19125 4031 19128
rect 3973 19119 4031 19125
rect 4614 19116 4620 19168
rect 4672 19116 4678 19168
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 6457 19159 6515 19165
rect 6457 19156 6469 19159
rect 6052 19128 6469 19156
rect 6052 19116 6058 19128
rect 6457 19125 6469 19128
rect 6503 19125 6515 19159
rect 6457 19119 6515 19125
rect 11330 19116 11336 19168
rect 11388 19116 11394 19168
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 12676 19128 13829 19156
rect 12676 19116 12682 19128
rect 13817 19125 13829 19128
rect 13863 19156 13875 19159
rect 14274 19156 14280 19168
rect 13863 19128 14280 19156
rect 13863 19125 13875 19128
rect 13817 19119 13875 19125
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 16224 19165 16252 19196
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 16669 19227 16727 19233
rect 16669 19193 16681 19227
rect 16715 19224 16727 19227
rect 17310 19224 17316 19236
rect 16715 19196 17316 19224
rect 16715 19193 16727 19196
rect 16669 19187 16727 19193
rect 17310 19184 17316 19196
rect 17368 19184 17374 19236
rect 17604 19224 17632 19264
rect 17957 19295 18015 19301
rect 17957 19261 17969 19295
rect 18003 19292 18015 19295
rect 18003 19264 18276 19292
rect 18003 19261 18015 19264
rect 17957 19255 18015 19261
rect 18248 19236 18276 19264
rect 18506 19252 18512 19304
rect 18564 19252 18570 19304
rect 20548 19292 20576 19323
rect 21082 19320 21088 19332
rect 21140 19360 21146 19372
rect 21468 19369 21496 19400
rect 21634 19388 21640 19440
rect 21692 19428 21698 19440
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 21692 19400 22385 19428
rect 21692 19388 21698 19400
rect 22373 19397 22385 19400
rect 22419 19397 22431 19431
rect 22373 19391 22431 19397
rect 21177 19363 21235 19369
rect 21177 19360 21189 19363
rect 21140 19332 21189 19360
rect 21140 19320 21146 19332
rect 21177 19329 21189 19332
rect 21223 19329 21235 19363
rect 21177 19323 21235 19329
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 21818 19320 21824 19372
rect 21876 19360 21882 19372
rect 21876 19332 21956 19360
rect 21876 19320 21882 19332
rect 20364 19264 20576 19292
rect 18138 19224 18144 19236
rect 17604 19196 18144 19224
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18230 19184 18236 19236
rect 18288 19184 18294 19236
rect 16209 19159 16267 19165
rect 16209 19125 16221 19159
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 17034 19116 17040 19168
rect 17092 19116 17098 19168
rect 17218 19116 17224 19168
rect 17276 19116 17282 19168
rect 17402 19116 17408 19168
rect 17460 19156 17466 19168
rect 19245 19159 19303 19165
rect 19245 19156 19257 19159
rect 17460 19128 19257 19156
rect 17460 19116 17466 19128
rect 19245 19125 19257 19128
rect 19291 19125 19303 19159
rect 19245 19119 19303 19125
rect 20073 19159 20131 19165
rect 20073 19125 20085 19159
rect 20119 19156 20131 19159
rect 20364 19156 20392 19264
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 21361 19295 21419 19301
rect 21361 19292 21373 19295
rect 20772 19264 21373 19292
rect 20772 19252 20778 19264
rect 21361 19261 21373 19264
rect 21407 19261 21419 19295
rect 21928 19292 21956 19332
rect 22002 19320 22008 19372
rect 22060 19320 22066 19372
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 22112 19332 22293 19360
rect 22112 19292 22140 19332
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 22281 19323 22339 19329
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19360 23167 19363
rect 23382 19360 23388 19372
rect 23155 19332 23388 19360
rect 23155 19329 23167 19332
rect 23109 19323 23167 19329
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 21928 19264 22140 19292
rect 21361 19255 21419 19261
rect 20438 19184 20444 19236
rect 20496 19224 20502 19236
rect 20625 19227 20683 19233
rect 20625 19224 20637 19227
rect 20496 19196 20637 19224
rect 20496 19184 20502 19196
rect 20625 19193 20637 19196
rect 20671 19193 20683 19227
rect 21269 19227 21327 19233
rect 21269 19224 21281 19227
rect 20625 19187 20683 19193
rect 20732 19196 21281 19224
rect 20732 19156 20760 19196
rect 21269 19193 21281 19196
rect 21315 19224 21327 19227
rect 21450 19224 21456 19236
rect 21315 19196 21456 19224
rect 21315 19193 21327 19196
rect 21269 19187 21327 19193
rect 21450 19184 21456 19196
rect 21508 19224 21514 19236
rect 22002 19224 22008 19236
rect 21508 19196 22008 19224
rect 21508 19184 21514 19196
rect 22002 19184 22008 19196
rect 22060 19184 22066 19236
rect 20119 19128 20760 19156
rect 20993 19159 21051 19165
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 20993 19125 21005 19159
rect 21039 19156 21051 19159
rect 21542 19156 21548 19168
rect 21039 19128 21548 19156
rect 21039 19125 21051 19128
rect 20993 19119 21051 19125
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 1104 19066 26312 19088
rect 1104 19014 4101 19066
rect 4153 19014 4165 19066
rect 4217 19014 4229 19066
rect 4281 19014 4293 19066
rect 4345 19014 4357 19066
rect 4409 19014 10403 19066
rect 10455 19014 10467 19066
rect 10519 19014 10531 19066
rect 10583 19014 10595 19066
rect 10647 19014 10659 19066
rect 10711 19014 16705 19066
rect 16757 19014 16769 19066
rect 16821 19014 16833 19066
rect 16885 19014 16897 19066
rect 16949 19014 16961 19066
rect 17013 19014 23007 19066
rect 23059 19014 23071 19066
rect 23123 19014 23135 19066
rect 23187 19014 23199 19066
rect 23251 19014 23263 19066
rect 23315 19014 26312 19066
rect 1104 18992 26312 19014
rect 2409 18955 2467 18961
rect 2409 18921 2421 18955
rect 2455 18952 2467 18955
rect 2774 18952 2780 18964
rect 2455 18924 2780 18952
rect 2455 18921 2467 18924
rect 2409 18915 2467 18921
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 6454 18912 6460 18964
rect 6512 18952 6518 18964
rect 6549 18955 6607 18961
rect 6549 18952 6561 18955
rect 6512 18924 6561 18952
rect 6512 18912 6518 18924
rect 6549 18921 6561 18924
rect 6595 18921 6607 18955
rect 6549 18915 6607 18921
rect 7190 18912 7196 18964
rect 7248 18912 7254 18964
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 9769 18955 9827 18961
rect 9769 18952 9781 18955
rect 9732 18924 9781 18952
rect 9732 18912 9738 18924
rect 9769 18921 9781 18924
rect 9815 18921 9827 18955
rect 9769 18915 9827 18921
rect 10965 18955 11023 18961
rect 10965 18921 10977 18955
rect 11011 18952 11023 18955
rect 11422 18952 11428 18964
rect 11011 18924 11428 18952
rect 11011 18921 11023 18924
rect 10965 18915 11023 18921
rect 11422 18912 11428 18924
rect 11480 18912 11486 18964
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 19242 18952 19248 18964
rect 14608 18924 19248 18952
rect 14608 18912 14614 18924
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19567 18955 19625 18961
rect 19567 18952 19579 18955
rect 19392 18924 19579 18952
rect 19392 18912 19398 18924
rect 19567 18921 19579 18924
rect 19613 18952 19625 18955
rect 20070 18952 20076 18964
rect 19613 18924 20076 18952
rect 19613 18921 19625 18924
rect 19567 18915 19625 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 20254 18912 20260 18964
rect 20312 18912 20318 18964
rect 20441 18955 20499 18961
rect 20441 18921 20453 18955
rect 20487 18952 20499 18955
rect 20622 18952 20628 18964
rect 20487 18924 20628 18952
rect 20487 18921 20499 18924
rect 20441 18915 20499 18921
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21082 18952 21088 18964
rect 20772 18924 21088 18952
rect 20772 18912 20778 18924
rect 21082 18912 21088 18924
rect 21140 18952 21146 18964
rect 23845 18955 23903 18961
rect 23845 18952 23857 18955
rect 21140 18924 23857 18952
rect 21140 18912 21146 18924
rect 23845 18921 23857 18924
rect 23891 18921 23903 18955
rect 23845 18915 23903 18921
rect 14458 18844 14464 18896
rect 14516 18844 14522 18896
rect 16393 18887 16451 18893
rect 16393 18853 16405 18887
rect 16439 18884 16451 18887
rect 16482 18884 16488 18896
rect 16439 18856 16488 18884
rect 16439 18853 16451 18856
rect 16393 18847 16451 18853
rect 16482 18844 16488 18856
rect 16540 18844 16546 18896
rect 17034 18844 17040 18896
rect 17092 18884 17098 18896
rect 20272 18884 20300 18912
rect 17092 18856 17632 18884
rect 17092 18844 17098 18856
rect 5258 18776 5264 18828
rect 5316 18816 5322 18828
rect 5534 18816 5540 18828
rect 5316 18788 5540 18816
rect 5316 18776 5322 18788
rect 5534 18776 5540 18788
rect 5592 18776 5598 18828
rect 6362 18776 6368 18828
rect 6420 18816 6426 18828
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 6420 18788 7389 18816
rect 6420 18776 6426 18788
rect 7377 18785 7389 18788
rect 7423 18785 7435 18819
rect 7377 18779 7435 18785
rect 10318 18776 10324 18828
rect 10376 18776 10382 18828
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 15749 18819 15807 18825
rect 13219 18788 14596 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 2314 18708 2320 18760
rect 2372 18708 2378 18760
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18748 5043 18751
rect 6546 18748 6552 18760
rect 5031 18720 6552 18748
rect 5031 18717 5043 18720
rect 4985 18711 5043 18717
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 7098 18708 7104 18760
rect 7156 18708 7162 18760
rect 10873 18751 10931 18757
rect 10873 18717 10885 18751
rect 10919 18748 10931 18751
rect 11514 18748 11520 18760
rect 10919 18720 11520 18748
rect 10919 18717 10931 18720
rect 10873 18711 10931 18717
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 12621 18751 12679 18757
rect 12621 18748 12633 18751
rect 12406 18720 12633 18748
rect 5258 18640 5264 18692
rect 5316 18640 5322 18692
rect 10229 18683 10287 18689
rect 10229 18649 10241 18683
rect 10275 18680 10287 18683
rect 11330 18680 11336 18692
rect 10275 18652 11336 18680
rect 10275 18649 10287 18652
rect 10229 18643 10287 18649
rect 11330 18640 11336 18652
rect 11388 18680 11394 18692
rect 12406 18680 12434 18720
rect 12621 18717 12633 18720
rect 12667 18748 12679 18751
rect 12986 18748 12992 18760
rect 12667 18720 12992 18748
rect 12667 18717 12679 18720
rect 12621 18711 12679 18717
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 13262 18708 13268 18760
rect 13320 18708 13326 18760
rect 14366 18748 14372 18760
rect 13556 18720 14372 18748
rect 11388 18652 12434 18680
rect 11388 18640 11394 18652
rect 12710 18640 12716 18692
rect 12768 18680 12774 18692
rect 13556 18689 13584 18720
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14568 18757 14596 18788
rect 15749 18785 15761 18819
rect 15795 18816 15807 18819
rect 15795 18788 17264 18816
rect 15795 18785 15807 18788
rect 15749 18779 15807 18785
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 15930 18708 15936 18760
rect 15988 18708 15994 18760
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 17236 18757 17264 18788
rect 16209 18751 16267 18757
rect 16209 18748 16221 18751
rect 16172 18720 16221 18748
rect 16172 18708 16178 18720
rect 16209 18717 16221 18720
rect 16255 18717 16267 18751
rect 16209 18711 16267 18717
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18717 17279 18751
rect 17221 18711 17279 18717
rect 17310 18708 17316 18760
rect 17368 18748 17374 18760
rect 17604 18757 17632 18856
rect 19444 18856 21220 18884
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 17368 18720 17509 18748
rect 17368 18708 17374 18720
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18748 17647 18751
rect 17770 18748 17776 18760
rect 17635 18720 17776 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18748 17923 18751
rect 17954 18748 17960 18760
rect 17911 18720 17960 18748
rect 17911 18717 17923 18720
rect 17865 18711 17923 18717
rect 17954 18708 17960 18720
rect 18012 18748 18018 18760
rect 19444 18757 19472 18856
rect 20070 18776 20076 18828
rect 20128 18816 20134 18828
rect 20128 18788 20944 18816
rect 20128 18776 20134 18788
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 18012 18720 18337 18748
rect 18012 18708 18018 18720
rect 18325 18717 18337 18720
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 18555 18720 19441 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 19705 18751 19763 18757
rect 19705 18748 19717 18751
rect 19668 18720 19717 18748
rect 19668 18708 19674 18720
rect 19705 18717 19717 18720
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 13541 18683 13599 18689
rect 13541 18680 13553 18683
rect 12768 18652 13553 18680
rect 12768 18640 12774 18652
rect 13541 18649 13553 18652
rect 13587 18649 13599 18683
rect 13541 18643 13599 18649
rect 13630 18640 13636 18692
rect 13688 18680 13694 18692
rect 14093 18683 14151 18689
rect 14093 18680 14105 18683
rect 13688 18652 14105 18680
rect 13688 18640 13694 18652
rect 14093 18649 14105 18652
rect 14139 18680 14151 18683
rect 14182 18680 14188 18692
rect 14139 18652 14188 18680
rect 14139 18649 14151 18652
rect 14093 18643 14151 18649
rect 14182 18640 14188 18652
rect 14240 18680 14246 18692
rect 14645 18683 14703 18689
rect 14645 18680 14657 18683
rect 14240 18652 14657 18680
rect 14240 18640 14246 18652
rect 14645 18649 14657 18652
rect 14691 18680 14703 18683
rect 14826 18680 14832 18692
rect 14691 18652 14832 18680
rect 14691 18649 14703 18652
rect 14645 18643 14703 18649
rect 14826 18640 14832 18652
rect 14884 18640 14890 18692
rect 16390 18640 16396 18692
rect 16448 18640 16454 18692
rect 17129 18683 17187 18689
rect 17129 18680 17141 18683
rect 16500 18652 17141 18680
rect 5077 18615 5135 18621
rect 5077 18581 5089 18615
rect 5123 18612 5135 18615
rect 5166 18612 5172 18624
rect 5123 18584 5172 18612
rect 5123 18581 5135 18584
rect 5077 18575 5135 18581
rect 5166 18572 5172 18584
rect 5224 18572 5230 18624
rect 7653 18615 7711 18621
rect 7653 18581 7665 18615
rect 7699 18612 7711 18615
rect 8754 18612 8760 18624
rect 7699 18584 8760 18612
rect 7699 18581 7711 18584
rect 7653 18575 7711 18581
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 10134 18572 10140 18624
rect 10192 18572 10198 18624
rect 12894 18572 12900 18624
rect 12952 18612 12958 18624
rect 14293 18615 14351 18621
rect 14293 18612 14305 18615
rect 12952 18584 14305 18612
rect 12952 18572 12958 18584
rect 14293 18581 14305 18584
rect 14339 18581 14351 18615
rect 14293 18575 14351 18581
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15804 18584 16129 18612
rect 15804 18572 15810 18584
rect 16117 18581 16129 18584
rect 16163 18612 16175 18615
rect 16500 18612 16528 18652
rect 17129 18649 17141 18652
rect 17175 18649 17187 18683
rect 17129 18643 17187 18649
rect 17405 18683 17463 18689
rect 17405 18649 17417 18683
rect 17451 18649 17463 18683
rect 17405 18643 17463 18649
rect 18049 18683 18107 18689
rect 18049 18649 18061 18683
rect 18095 18680 18107 18683
rect 19720 18680 19748 18711
rect 19794 18708 19800 18760
rect 19852 18748 19858 18760
rect 19889 18751 19947 18757
rect 19889 18748 19901 18751
rect 19852 18720 19901 18748
rect 19852 18708 19858 18720
rect 19889 18717 19901 18720
rect 19935 18748 19947 18751
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 19935 18720 20269 18748
rect 19935 18717 19947 18720
rect 19889 18711 19947 18717
rect 20257 18717 20269 18720
rect 20303 18748 20315 18751
rect 20714 18748 20720 18760
rect 20303 18720 20720 18748
rect 20303 18717 20315 18720
rect 20257 18711 20315 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 20916 18757 20944 18788
rect 21082 18776 21088 18828
rect 21140 18776 21146 18828
rect 20809 18751 20867 18757
rect 20809 18717 20821 18751
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 20993 18751 21051 18757
rect 20993 18717 21005 18751
rect 21039 18748 21051 18751
rect 21192 18748 21220 18856
rect 23474 18844 23480 18896
rect 23532 18884 23538 18896
rect 23532 18856 23980 18884
rect 23532 18844 23538 18856
rect 21039 18720 21220 18748
rect 21039 18717 21051 18720
rect 20993 18711 21051 18717
rect 19981 18683 20039 18689
rect 19981 18680 19993 18683
rect 18095 18652 19334 18680
rect 19720 18652 19993 18680
rect 18095 18649 18107 18652
rect 18049 18643 18107 18649
rect 16163 18584 16528 18612
rect 16163 18581 16175 18584
rect 16117 18575 16175 18581
rect 16850 18572 16856 18624
rect 16908 18572 16914 18624
rect 16945 18615 17003 18621
rect 16945 18581 16957 18615
rect 16991 18612 17003 18615
rect 17034 18612 17040 18624
rect 16991 18584 17040 18612
rect 16991 18581 17003 18584
rect 16945 18575 17003 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 17420 18612 17448 18643
rect 17276 18584 17448 18612
rect 17276 18572 17282 18584
rect 17770 18572 17776 18624
rect 17828 18572 17834 18624
rect 18230 18572 18236 18624
rect 18288 18572 18294 18624
rect 18690 18572 18696 18624
rect 18748 18572 18754 18624
rect 19306 18612 19334 18652
rect 19981 18649 19993 18652
rect 20027 18649 20039 18683
rect 19981 18643 20039 18649
rect 20530 18640 20536 18692
rect 20588 18680 20594 18692
rect 20824 18680 20852 18711
rect 21266 18708 21272 18760
rect 21324 18708 21330 18760
rect 21358 18708 21364 18760
rect 21416 18748 21422 18760
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 21416 18720 21649 18748
rect 21416 18708 21422 18720
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 22094 18708 22100 18760
rect 22152 18708 22158 18760
rect 23952 18757 23980 18856
rect 23937 18751 23995 18757
rect 23937 18717 23949 18751
rect 23983 18717 23995 18751
rect 23937 18711 23995 18717
rect 20588 18652 20852 18680
rect 20588 18640 20594 18652
rect 21450 18640 21456 18692
rect 21508 18640 21514 18692
rect 21542 18640 21548 18692
rect 21600 18640 21606 18692
rect 22373 18683 22431 18689
rect 22373 18680 22385 18683
rect 22066 18652 22385 18680
rect 19794 18612 19800 18624
rect 19306 18584 19800 18612
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 19889 18615 19947 18621
rect 19889 18581 19901 18615
rect 19935 18612 19947 18615
rect 20346 18612 20352 18624
rect 19935 18584 20352 18612
rect 19935 18581 19947 18584
rect 19889 18575 19947 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 20625 18615 20683 18621
rect 20625 18581 20637 18615
rect 20671 18612 20683 18615
rect 21082 18612 21088 18624
rect 20671 18584 21088 18612
rect 20671 18581 20683 18584
rect 20625 18575 20683 18581
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 21821 18615 21879 18621
rect 21821 18581 21833 18615
rect 21867 18612 21879 18615
rect 22066 18612 22094 18652
rect 22373 18649 22385 18652
rect 22419 18649 22431 18683
rect 24029 18683 24087 18689
rect 24029 18680 24041 18683
rect 23598 18652 24041 18680
rect 22373 18643 22431 18649
rect 24029 18649 24041 18652
rect 24075 18649 24087 18683
rect 24029 18643 24087 18649
rect 21867 18584 22094 18612
rect 21867 18581 21879 18584
rect 21821 18575 21879 18581
rect 1104 18522 26312 18544
rect 1104 18470 4761 18522
rect 4813 18470 4825 18522
rect 4877 18470 4889 18522
rect 4941 18470 4953 18522
rect 5005 18470 5017 18522
rect 5069 18470 11063 18522
rect 11115 18470 11127 18522
rect 11179 18470 11191 18522
rect 11243 18470 11255 18522
rect 11307 18470 11319 18522
rect 11371 18470 17365 18522
rect 17417 18470 17429 18522
rect 17481 18470 17493 18522
rect 17545 18470 17557 18522
rect 17609 18470 17621 18522
rect 17673 18470 23667 18522
rect 23719 18470 23731 18522
rect 23783 18470 23795 18522
rect 23847 18470 23859 18522
rect 23911 18470 23923 18522
rect 23975 18470 26312 18522
rect 1104 18448 26312 18470
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18377 2651 18411
rect 2593 18371 2651 18377
rect 2961 18411 3019 18417
rect 2961 18377 2973 18411
rect 3007 18408 3019 18411
rect 3786 18408 3792 18420
rect 3007 18380 3792 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2608 18272 2636 18371
rect 3786 18368 3792 18380
rect 3844 18408 3850 18420
rect 4249 18411 4307 18417
rect 4249 18408 4261 18411
rect 3844 18380 4261 18408
rect 3844 18368 3850 18380
rect 4249 18377 4261 18380
rect 4295 18377 4307 18411
rect 4249 18371 4307 18377
rect 5258 18368 5264 18420
rect 5316 18408 5322 18420
rect 7653 18411 7711 18417
rect 7653 18408 7665 18411
rect 5316 18380 7665 18408
rect 5316 18368 5322 18380
rect 7653 18377 7665 18380
rect 7699 18377 7711 18411
rect 7653 18371 7711 18377
rect 8570 18368 8576 18420
rect 8628 18368 8634 18420
rect 10778 18408 10784 18420
rect 9646 18380 10784 18408
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 6365 18343 6423 18349
rect 6365 18340 6377 18343
rect 3292 18312 6377 18340
rect 3292 18300 3298 18312
rect 6365 18309 6377 18312
rect 6411 18309 6423 18343
rect 6365 18303 6423 18309
rect 8665 18343 8723 18349
rect 8665 18309 8677 18343
rect 8711 18340 8723 18343
rect 9306 18340 9312 18352
rect 8711 18312 9312 18340
rect 8711 18309 8723 18312
rect 8665 18303 8723 18309
rect 9306 18300 9312 18312
rect 9364 18300 9370 18352
rect 2363 18244 2636 18272
rect 3789 18275 3847 18281
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 3789 18241 3801 18275
rect 3835 18272 3847 18275
rect 4341 18275 4399 18281
rect 3835 18244 3924 18272
rect 3835 18241 3847 18244
rect 3789 18235 3847 18241
rect 3050 18164 3056 18216
rect 3108 18164 3114 18216
rect 3237 18207 3295 18213
rect 3237 18173 3249 18207
rect 3283 18204 3295 18207
rect 3602 18204 3608 18216
rect 3283 18176 3608 18204
rect 3283 18173 3295 18176
rect 3237 18167 3295 18173
rect 3602 18164 3608 18176
rect 3660 18164 3666 18216
rect 3896 18145 3924 18244
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 4387 18244 4660 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 4430 18164 4436 18216
rect 4488 18164 4494 18216
rect 4632 18204 4660 18244
rect 4706 18232 4712 18284
rect 4764 18232 4770 18284
rect 4908 18244 5212 18272
rect 4908 18204 4936 18244
rect 4632 18176 4936 18204
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18204 5043 18207
rect 5074 18204 5080 18216
rect 5031 18176 5080 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5184 18204 5212 18244
rect 5350 18232 5356 18284
rect 5408 18272 5414 18284
rect 5813 18275 5871 18281
rect 5813 18272 5825 18275
rect 5408 18244 5825 18272
rect 5408 18232 5414 18244
rect 5813 18241 5825 18244
rect 5859 18241 5871 18275
rect 5813 18235 5871 18241
rect 5184 18176 5396 18204
rect 3881 18139 3939 18145
rect 3881 18105 3893 18139
rect 3927 18105 3939 18139
rect 3881 18099 3939 18105
rect 4522 18096 4528 18148
rect 4580 18136 4586 18148
rect 5261 18139 5319 18145
rect 5261 18136 5273 18139
rect 4580 18108 5273 18136
rect 4580 18096 4586 18108
rect 5261 18105 5273 18108
rect 5307 18105 5319 18139
rect 5368 18136 5396 18176
rect 5442 18164 5448 18216
rect 5500 18164 5506 18216
rect 5828 18204 5856 18235
rect 5994 18232 6000 18284
rect 6052 18232 6058 18284
rect 6178 18232 6184 18284
rect 6236 18232 6242 18284
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18241 9275 18275
rect 9324 18272 9352 18300
rect 9646 18272 9674 18380
rect 10778 18368 10784 18380
rect 10836 18408 10842 18420
rect 11882 18408 11888 18420
rect 10836 18380 11888 18408
rect 10836 18368 10842 18380
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 14093 18411 14151 18417
rect 14093 18377 14105 18411
rect 14139 18408 14151 18411
rect 14550 18408 14556 18420
rect 14139 18380 14556 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 10318 18300 10324 18352
rect 10376 18340 10382 18352
rect 10689 18343 10747 18349
rect 10689 18340 10701 18343
rect 10376 18312 10701 18340
rect 10376 18300 10382 18312
rect 10689 18309 10701 18312
rect 10735 18340 10747 18343
rect 10735 18312 12388 18340
rect 10735 18309 10747 18312
rect 10689 18303 10747 18309
rect 9324 18244 9674 18272
rect 10597 18275 10655 18281
rect 9217 18235 9275 18241
rect 10597 18241 10609 18275
rect 10643 18241 10655 18275
rect 10597 18235 10655 18241
rect 6822 18204 6828 18216
rect 5828 18176 6828 18204
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 8754 18164 8760 18216
rect 8812 18164 8818 18216
rect 5626 18136 5632 18148
rect 5368 18108 5632 18136
rect 5261 18099 5319 18105
rect 5626 18096 5632 18108
rect 5684 18096 5690 18148
rect 8205 18139 8263 18145
rect 8205 18105 8217 18139
rect 8251 18136 8263 18139
rect 9232 18136 9260 18235
rect 9950 18164 9956 18216
rect 10008 18204 10014 18216
rect 10618 18204 10646 18235
rect 10778 18232 10784 18284
rect 10836 18232 10842 18284
rect 10870 18232 10876 18284
rect 10928 18232 10934 18284
rect 11054 18232 11060 18284
rect 11112 18232 11118 18284
rect 11164 18244 11652 18272
rect 11164 18204 11192 18244
rect 10008 18176 11192 18204
rect 11241 18207 11299 18213
rect 10008 18164 10014 18176
rect 11241 18173 11253 18207
rect 11287 18204 11299 18207
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 11287 18176 11529 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 11624 18204 11652 18244
rect 11698 18232 11704 18284
rect 11756 18232 11762 18284
rect 11882 18232 11888 18284
rect 11940 18232 11946 18284
rect 12360 18281 12388 18312
rect 12912 18312 13676 18340
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12618 18232 12624 18284
rect 12676 18272 12682 18284
rect 12912 18281 12940 18312
rect 12897 18275 12955 18281
rect 12897 18272 12909 18275
rect 12676 18244 12909 18272
rect 12676 18232 12682 18244
rect 12897 18241 12909 18244
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 13538 18232 13544 18284
rect 13596 18232 13602 18284
rect 13648 18281 13676 18312
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18241 13691 18275
rect 13633 18235 13691 18241
rect 13906 18232 13912 18284
rect 13964 18232 13970 18284
rect 11790 18204 11796 18216
rect 11624 18176 11796 18204
rect 11517 18167 11575 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 11977 18207 12035 18213
rect 11977 18173 11989 18207
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 12161 18207 12219 18213
rect 12161 18173 12173 18207
rect 12207 18204 12219 18207
rect 14108 18204 14136 18371
rect 14550 18368 14556 18380
rect 14608 18368 14614 18420
rect 15930 18368 15936 18420
rect 15988 18408 15994 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 15988 18380 16681 18408
rect 15988 18368 15994 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 16669 18371 16727 18377
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 17589 18411 17647 18417
rect 17589 18408 17601 18411
rect 17000 18380 17601 18408
rect 17000 18368 17006 18380
rect 17589 18377 17601 18380
rect 17635 18377 17647 18411
rect 17589 18371 17647 18377
rect 17954 18368 17960 18420
rect 18012 18417 18018 18420
rect 18012 18411 18041 18417
rect 18029 18408 18041 18411
rect 18690 18408 18696 18420
rect 18029 18380 18696 18408
rect 18029 18377 18041 18380
rect 18012 18371 18041 18377
rect 18012 18368 18018 18371
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 19702 18368 19708 18420
rect 19760 18408 19766 18420
rect 19997 18411 20055 18417
rect 19997 18408 20009 18411
rect 19760 18380 20009 18408
rect 19760 18368 19766 18380
rect 19997 18377 20009 18380
rect 20043 18377 20055 18411
rect 19997 18371 20055 18377
rect 20162 18368 20168 18420
rect 20220 18368 20226 18420
rect 20625 18411 20683 18417
rect 20625 18377 20637 18411
rect 20671 18408 20683 18411
rect 20671 18380 21312 18408
rect 20671 18377 20683 18380
rect 20625 18371 20683 18377
rect 16114 18300 16120 18352
rect 16172 18300 16178 18352
rect 16333 18343 16391 18349
rect 16333 18309 16345 18343
rect 16379 18340 16391 18343
rect 17773 18343 17831 18349
rect 16379 18312 17372 18340
rect 16379 18309 16391 18312
rect 16333 18303 16391 18309
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18272 14427 18275
rect 14642 18272 14648 18284
rect 14415 18244 14648 18272
rect 14415 18241 14427 18244
rect 14369 18235 14427 18241
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 14826 18232 14832 18284
rect 14884 18232 14890 18284
rect 16850 18232 16856 18284
rect 16908 18272 16914 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16908 18244 17233 18272
rect 16908 18232 16914 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 12207 18176 14136 18204
rect 14185 18207 14243 18213
rect 12207 18173 12219 18176
rect 12161 18167 12219 18173
rect 14185 18173 14197 18207
rect 14231 18173 14243 18207
rect 14185 18167 14243 18173
rect 17129 18207 17187 18213
rect 17129 18173 17141 18207
rect 17175 18173 17187 18207
rect 17344 18204 17372 18312
rect 17773 18309 17785 18343
rect 17819 18340 17831 18343
rect 18138 18340 18144 18352
rect 17819 18312 18144 18340
rect 17819 18309 17831 18312
rect 17773 18303 17831 18309
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 19794 18300 19800 18352
rect 19852 18300 19858 18352
rect 20346 18300 20352 18352
rect 20404 18340 20410 18352
rect 21284 18340 21312 18380
rect 21358 18368 21364 18420
rect 21416 18368 21422 18420
rect 25130 18368 25136 18420
rect 25188 18368 25194 18420
rect 21450 18340 21456 18352
rect 20404 18312 21220 18340
rect 21284 18312 21456 18340
rect 20404 18300 20410 18312
rect 17402 18232 17408 18284
rect 17460 18232 17466 18284
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18272 17739 18275
rect 18230 18272 18236 18284
rect 17727 18244 18236 18272
rect 17727 18241 17739 18244
rect 17681 18235 17739 18241
rect 17696 18204 17724 18235
rect 18230 18232 18236 18244
rect 18288 18232 18294 18284
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20772 18244 20821 18272
rect 20772 18232 20778 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20990 18232 20996 18284
rect 21048 18232 21054 18284
rect 21082 18232 21088 18284
rect 21140 18232 21146 18284
rect 21192 18281 21220 18312
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 21177 18275 21235 18281
rect 21177 18241 21189 18275
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 21361 18275 21419 18281
rect 21361 18241 21373 18275
rect 21407 18241 21419 18275
rect 21361 18235 21419 18241
rect 17344 18176 17724 18204
rect 17129 18167 17187 18173
rect 8251 18108 9260 18136
rect 11149 18139 11207 18145
rect 8251 18105 8263 18108
rect 8205 18099 8263 18105
rect 11149 18105 11161 18139
rect 11195 18136 11207 18139
rect 11992 18136 12020 18167
rect 12529 18139 12587 18145
rect 12529 18136 12541 18139
rect 11195 18108 11836 18136
rect 11992 18108 12541 18136
rect 11195 18105 11207 18108
rect 11149 18099 11207 18105
rect 1670 18028 1676 18080
rect 1728 18068 1734 18080
rect 2133 18071 2191 18077
rect 2133 18068 2145 18071
rect 1728 18040 2145 18068
rect 1728 18028 1734 18040
rect 2133 18037 2145 18040
rect 2179 18037 2191 18071
rect 2133 18031 2191 18037
rect 3602 18028 3608 18080
rect 3660 18028 3666 18080
rect 4798 18028 4804 18080
rect 4856 18028 4862 18080
rect 5350 18028 5356 18080
rect 5408 18028 5414 18080
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 5721 18071 5779 18077
rect 5721 18068 5733 18071
rect 5500 18040 5733 18068
rect 5500 18028 5506 18040
rect 5721 18037 5733 18040
rect 5767 18037 5779 18071
rect 5721 18031 5779 18037
rect 9030 18028 9036 18080
rect 9088 18028 9094 18080
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 10836 18040 11253 18068
rect 10836 18028 10842 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 11241 18031 11299 18037
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 11698 18068 11704 18080
rect 11388 18040 11704 18068
rect 11388 18028 11394 18040
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 11808 18068 11836 18108
rect 12529 18105 12541 18108
rect 12575 18105 12587 18139
rect 13078 18136 13084 18148
rect 12529 18099 12587 18105
rect 12912 18108 13084 18136
rect 12912 18068 12940 18108
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 14200 18136 14228 18167
rect 13280 18108 14228 18136
rect 11808 18040 12940 18068
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 13173 18071 13231 18077
rect 13173 18068 13185 18071
rect 13044 18040 13185 18068
rect 13044 18028 13050 18040
rect 13173 18037 13185 18040
rect 13219 18068 13231 18071
rect 13280 18068 13308 18108
rect 16482 18096 16488 18148
rect 16540 18136 16546 18148
rect 17144 18136 17172 18167
rect 20622 18164 20628 18216
rect 20680 18204 20686 18216
rect 21376 18204 21404 18235
rect 25038 18232 25044 18284
rect 25096 18232 25102 18284
rect 20680 18176 21404 18204
rect 20680 18164 20686 18176
rect 16540 18108 17172 18136
rect 16540 18096 16546 18108
rect 17218 18096 17224 18148
rect 17276 18096 17282 18148
rect 18141 18139 18199 18145
rect 18141 18136 18153 18139
rect 17328 18108 18153 18136
rect 13219 18040 13308 18068
rect 13219 18037 13231 18040
rect 13173 18031 13231 18037
rect 13354 18028 13360 18080
rect 13412 18028 13418 18080
rect 13814 18028 13820 18080
rect 13872 18028 13878 18080
rect 14550 18028 14556 18080
rect 14608 18028 14614 18080
rect 14737 18071 14795 18077
rect 14737 18037 14749 18071
rect 14783 18068 14795 18071
rect 15010 18068 15016 18080
rect 14783 18040 15016 18068
rect 14783 18037 14795 18040
rect 14737 18031 14795 18037
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 16206 18028 16212 18080
rect 16264 18068 16270 18080
rect 16301 18071 16359 18077
rect 16301 18068 16313 18071
rect 16264 18040 16313 18068
rect 16264 18028 16270 18040
rect 16301 18037 16313 18040
rect 16347 18068 16359 18071
rect 16942 18068 16948 18080
rect 16347 18040 16948 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 17236 18068 17264 18096
rect 17328 18068 17356 18108
rect 18141 18105 18153 18108
rect 18187 18105 18199 18139
rect 18141 18099 18199 18105
rect 20438 18096 20444 18148
rect 20496 18136 20502 18148
rect 20990 18136 20996 18148
rect 20496 18108 20996 18136
rect 20496 18096 20502 18108
rect 20990 18096 20996 18108
rect 21048 18096 21054 18148
rect 17083 18040 17356 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 17402 18028 17408 18080
rect 17460 18068 17466 18080
rect 17957 18071 18015 18077
rect 17957 18068 17969 18071
rect 17460 18040 17969 18068
rect 17460 18028 17466 18040
rect 17957 18037 17969 18040
rect 18003 18037 18015 18071
rect 17957 18031 18015 18037
rect 19794 18028 19800 18080
rect 19852 18068 19858 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19852 18040 19993 18068
rect 19852 18028 19858 18040
rect 19981 18037 19993 18040
rect 20027 18068 20039 18071
rect 20254 18068 20260 18080
rect 20027 18040 20260 18068
rect 20027 18037 20039 18040
rect 19981 18031 20039 18037
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 1104 17978 26312 18000
rect 1104 17926 4101 17978
rect 4153 17926 4165 17978
rect 4217 17926 4229 17978
rect 4281 17926 4293 17978
rect 4345 17926 4357 17978
rect 4409 17926 10403 17978
rect 10455 17926 10467 17978
rect 10519 17926 10531 17978
rect 10583 17926 10595 17978
rect 10647 17926 10659 17978
rect 10711 17926 16705 17978
rect 16757 17926 16769 17978
rect 16821 17926 16833 17978
rect 16885 17926 16897 17978
rect 16949 17926 16961 17978
rect 17013 17926 23007 17978
rect 23059 17926 23071 17978
rect 23123 17926 23135 17978
rect 23187 17926 23199 17978
rect 23251 17926 23263 17978
rect 23315 17926 26312 17978
rect 1104 17904 26312 17926
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 4856 17836 5166 17864
rect 4856 17824 4862 17836
rect 5138 17796 5166 17836
rect 5718 17824 5724 17876
rect 5776 17864 5782 17876
rect 6089 17867 6147 17873
rect 6089 17864 6101 17867
rect 5776 17836 6101 17864
rect 5776 17824 5782 17836
rect 6089 17833 6101 17836
rect 6135 17864 6147 17867
rect 6454 17864 6460 17876
rect 6135 17836 6460 17864
rect 6135 17833 6147 17836
rect 6089 17827 6147 17833
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 6730 17824 6736 17876
rect 6788 17864 6794 17876
rect 6917 17867 6975 17873
rect 6917 17864 6929 17867
rect 6788 17836 6929 17864
rect 6788 17824 6794 17836
rect 6917 17833 6929 17836
rect 6963 17833 6975 17867
rect 6917 17827 6975 17833
rect 7466 17824 7472 17876
rect 7524 17864 7530 17876
rect 13081 17867 13139 17873
rect 7524 17836 13032 17864
rect 7524 17824 7530 17836
rect 6178 17796 6184 17808
rect 5138 17768 6184 17796
rect 6178 17756 6184 17768
rect 6236 17796 6242 17808
rect 6748 17796 6776 17824
rect 6236 17768 6776 17796
rect 6236 17756 6242 17768
rect 7374 17756 7380 17808
rect 7432 17756 7438 17808
rect 7561 17799 7619 17805
rect 7561 17765 7573 17799
rect 7607 17796 7619 17799
rect 8386 17796 8392 17808
rect 7607 17768 8392 17796
rect 7607 17765 7619 17768
rect 7561 17759 7619 17765
rect 8386 17756 8392 17768
rect 8444 17756 8450 17808
rect 10226 17756 10232 17808
rect 10284 17796 10290 17808
rect 10870 17796 10876 17808
rect 10284 17768 10876 17796
rect 10284 17756 10290 17768
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 11882 17756 11888 17808
rect 11940 17796 11946 17808
rect 12529 17799 12587 17805
rect 12529 17796 12541 17799
rect 11940 17768 12541 17796
rect 11940 17756 11946 17768
rect 12529 17765 12541 17768
rect 12575 17765 12587 17799
rect 12529 17759 12587 17765
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 1412 17700 3801 17728
rect 1412 17672 1440 17700
rect 3789 17697 3801 17700
rect 3835 17728 3847 17731
rect 4430 17728 4436 17740
rect 3835 17700 4436 17728
rect 3835 17697 3847 17700
rect 3789 17691 3847 17697
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 5074 17688 5080 17740
rect 5132 17728 5138 17740
rect 5534 17728 5540 17740
rect 5132 17700 5540 17728
rect 5132 17688 5138 17700
rect 5534 17688 5540 17700
rect 5592 17728 5598 17740
rect 6733 17731 6791 17737
rect 5592 17700 5856 17728
rect 5592 17688 5598 17700
rect 1394 17620 1400 17672
rect 1452 17620 1458 17672
rect 3050 17620 3056 17672
rect 3108 17660 3114 17672
rect 3326 17660 3332 17672
rect 3108 17632 3332 17660
rect 3108 17620 3114 17632
rect 3326 17620 3332 17632
rect 3384 17660 3390 17672
rect 3421 17663 3479 17669
rect 3421 17660 3433 17663
rect 3384 17632 3433 17660
rect 3384 17620 3390 17632
rect 3421 17629 3433 17632
rect 3467 17629 3479 17663
rect 3421 17623 3479 17629
rect 5166 17620 5172 17672
rect 5224 17620 5230 17672
rect 5350 17620 5356 17672
rect 5408 17660 5414 17672
rect 5721 17663 5779 17669
rect 5721 17660 5733 17663
rect 5408 17632 5733 17660
rect 5408 17620 5414 17632
rect 1670 17552 1676 17604
rect 1728 17552 1734 17604
rect 2406 17552 2412 17604
rect 2464 17552 2470 17604
rect 3602 17552 3608 17604
rect 3660 17592 3666 17604
rect 4065 17595 4123 17601
rect 4065 17592 4077 17595
rect 3660 17564 4077 17592
rect 3660 17552 3666 17564
rect 4065 17561 4077 17564
rect 4111 17561 4123 17595
rect 4065 17555 4123 17561
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 5460 17524 5488 17632
rect 5721 17629 5733 17632
rect 5767 17629 5779 17663
rect 5721 17623 5779 17629
rect 5828 17592 5856 17700
rect 6733 17697 6745 17731
rect 6779 17728 6791 17731
rect 8113 17731 8171 17737
rect 8113 17728 8125 17731
rect 6779 17700 8125 17728
rect 6779 17697 6791 17700
rect 6733 17691 6791 17697
rect 8113 17697 8125 17700
rect 8159 17697 8171 17731
rect 8113 17691 8171 17697
rect 12066 17688 12072 17740
rect 12124 17688 12130 17740
rect 13004 17728 13032 17836
rect 13081 17833 13093 17867
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 13096 17796 13124 17827
rect 13170 17824 13176 17876
rect 13228 17864 13234 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 13228 17836 13277 17864
rect 13228 17824 13234 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13265 17827 13323 17833
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 13906 17864 13912 17876
rect 13771 17836 13912 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 14274 17824 14280 17876
rect 14332 17824 14338 17876
rect 16853 17867 16911 17873
rect 16853 17833 16865 17867
rect 16899 17864 16911 17867
rect 17034 17864 17040 17876
rect 16899 17836 17040 17864
rect 16899 17833 16911 17836
rect 16853 17827 16911 17833
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 13814 17796 13820 17808
rect 13096 17768 13820 17796
rect 13814 17756 13820 17768
rect 13872 17756 13878 17808
rect 18138 17796 18144 17808
rect 17052 17768 18144 17796
rect 16114 17728 16120 17740
rect 13004 17700 16120 17728
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6052 17632 6592 17660
rect 6052 17620 6058 17632
rect 6564 17601 6592 17632
rect 6638 17620 6644 17672
rect 6696 17660 6702 17672
rect 6822 17660 6828 17672
rect 6696 17632 6828 17660
rect 6696 17620 6702 17632
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 7098 17620 7104 17672
rect 7156 17620 7162 17672
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 7208 17632 8585 17660
rect 6365 17595 6423 17601
rect 6365 17592 6377 17595
rect 5828 17564 6377 17592
rect 6365 17561 6377 17564
rect 6411 17561 6423 17595
rect 6365 17555 6423 17561
rect 6549 17595 6607 17601
rect 6549 17561 6561 17595
rect 6595 17592 6607 17595
rect 7208 17592 7236 17632
rect 8573 17629 8585 17632
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17660 8999 17663
rect 9122 17660 9128 17672
rect 8987 17632 9128 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 10413 17663 10471 17669
rect 9999 17632 10364 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 6595 17564 7236 17592
rect 6595 17561 6607 17564
rect 6549 17555 6607 17561
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 8389 17595 8447 17601
rect 8389 17592 8401 17595
rect 7340 17564 8401 17592
rect 7340 17552 7346 17564
rect 8389 17561 8401 17564
rect 8435 17561 8447 17595
rect 8389 17555 8447 17561
rect 10134 17552 10140 17604
rect 10192 17552 10198 17604
rect 10336 17592 10364 17632
rect 10413 17629 10425 17663
rect 10459 17660 10471 17663
rect 12434 17660 12440 17672
rect 10459 17632 12440 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 12434 17620 12440 17632
rect 12492 17660 12498 17672
rect 13722 17660 13728 17672
rect 12492 17632 13728 17660
rect 12492 17620 12498 17632
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 17052 17669 17080 17768
rect 18138 17756 18144 17768
rect 18196 17756 18202 17808
rect 17954 17728 17960 17740
rect 17328 17700 17960 17728
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 14476 17632 14565 17660
rect 11514 17592 11520 17604
rect 10336 17564 11520 17592
rect 11514 17552 11520 17564
rect 11572 17552 11578 17604
rect 11790 17552 11796 17604
rect 11848 17592 11854 17604
rect 12253 17595 12311 17601
rect 12253 17592 12265 17595
rect 11848 17564 12265 17592
rect 11848 17552 11854 17564
rect 12253 17561 12265 17564
rect 12299 17561 12311 17595
rect 12253 17555 12311 17561
rect 12894 17552 12900 17604
rect 12952 17552 12958 17604
rect 13354 17552 13360 17604
rect 13412 17552 13418 17604
rect 13538 17552 13544 17604
rect 13596 17552 13602 17604
rect 14093 17595 14151 17601
rect 14093 17561 14105 17595
rect 14139 17592 14151 17595
rect 14182 17592 14188 17604
rect 14139 17564 14188 17592
rect 14139 17561 14151 17564
rect 14093 17555 14151 17561
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 4764 17496 5488 17524
rect 5537 17527 5595 17533
rect 4764 17484 4770 17496
rect 5537 17493 5549 17527
rect 5583 17524 5595 17527
rect 5626 17524 5632 17536
rect 5583 17496 5632 17524
rect 5583 17493 5595 17496
rect 5537 17487 5595 17493
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 6089 17527 6147 17533
rect 6089 17524 6101 17527
rect 6052 17496 6101 17524
rect 6052 17484 6058 17496
rect 6089 17493 6101 17496
rect 6135 17524 6147 17527
rect 6178 17524 6184 17536
rect 6135 17496 6184 17524
rect 6135 17493 6147 17496
rect 6089 17487 6147 17493
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 6270 17484 6276 17536
rect 6328 17484 6334 17536
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 7926 17524 7932 17536
rect 6696 17496 7932 17524
rect 6696 17484 6702 17496
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 8021 17527 8079 17533
rect 8021 17493 8033 17527
rect 8067 17524 8079 17527
rect 8662 17524 8668 17536
rect 8067 17496 8668 17524
rect 8067 17493 8079 17496
rect 8021 17487 8079 17493
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 8754 17484 8760 17536
rect 8812 17484 8818 17536
rect 8938 17484 8944 17536
rect 8996 17524 9002 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8996 17496 9045 17524
rect 8996 17484 9002 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 9033 17487 9091 17493
rect 10321 17527 10379 17533
rect 10321 17493 10333 17527
rect 10367 17524 10379 17527
rect 11422 17524 11428 17536
rect 10367 17496 11428 17524
rect 10367 17493 10379 17496
rect 10321 17487 10379 17493
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 12713 17527 12771 17533
rect 12713 17524 12725 17527
rect 12584 17496 12725 17524
rect 12584 17484 12590 17496
rect 12713 17493 12725 17496
rect 12759 17524 12771 17527
rect 13097 17527 13155 17533
rect 13097 17524 13109 17527
rect 12759 17496 13109 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 13097 17493 13109 17496
rect 13143 17493 13155 17527
rect 13097 17487 13155 17493
rect 13906 17484 13912 17536
rect 13964 17524 13970 17536
rect 14476 17533 14504 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 14553 17623 14611 17629
rect 17037 17663 17095 17669
rect 17037 17629 17049 17663
rect 17083 17629 17095 17663
rect 17037 17623 17095 17629
rect 17126 17620 17132 17672
rect 17184 17660 17190 17672
rect 17328 17669 17356 17700
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 19521 17731 19579 17737
rect 19521 17697 19533 17731
rect 19567 17728 19579 17731
rect 20070 17728 20076 17740
rect 19567 17700 20076 17728
rect 19567 17697 19579 17700
rect 19521 17691 19579 17697
rect 20070 17688 20076 17700
rect 20128 17728 20134 17740
rect 20254 17728 20260 17740
rect 20128 17700 20260 17728
rect 20128 17688 20134 17700
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 23474 17728 23480 17740
rect 22664 17700 23480 17728
rect 17221 17663 17279 17669
rect 17221 17660 17233 17663
rect 17184 17632 17233 17660
rect 17184 17620 17190 17632
rect 17221 17629 17233 17632
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17629 17555 17663
rect 19610 17660 19616 17672
rect 17497 17623 17555 17629
rect 18432 17632 19616 17660
rect 14293 17527 14351 17533
rect 14293 17524 14305 17527
rect 13964 17496 14305 17524
rect 13964 17484 13970 17496
rect 14293 17493 14305 17496
rect 14339 17493 14351 17527
rect 14293 17487 14351 17493
rect 14461 17527 14519 17533
rect 14461 17493 14473 17527
rect 14507 17493 14519 17527
rect 14461 17487 14519 17493
rect 14734 17484 14740 17536
rect 14792 17484 14798 17536
rect 14826 17484 14832 17536
rect 14884 17524 14890 17536
rect 17512 17524 17540 17623
rect 18141 17595 18199 17601
rect 18141 17561 18153 17595
rect 18187 17592 18199 17595
rect 18230 17592 18236 17604
rect 18187 17564 18236 17592
rect 18187 17561 18199 17564
rect 18141 17555 18199 17561
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 18432 17536 18460 17632
rect 19610 17620 19616 17632
rect 19668 17660 19674 17672
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19668 17632 19717 17660
rect 19668 17620 19674 17632
rect 19705 17629 19717 17632
rect 19751 17660 19763 17663
rect 19886 17660 19892 17672
rect 19751 17632 19892 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 19886 17620 19892 17632
rect 19944 17660 19950 17672
rect 20530 17660 20536 17672
rect 19944 17632 20536 17660
rect 19944 17620 19950 17632
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17660 21143 17663
rect 21174 17660 21180 17672
rect 21131 17632 21180 17660
rect 21131 17629 21143 17632
rect 21085 17623 21143 17629
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 21450 17620 21456 17672
rect 21508 17620 21514 17672
rect 22664 17669 22692 17700
rect 23474 17688 23480 17700
rect 23532 17688 23538 17740
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 23201 17663 23259 17669
rect 23201 17629 23213 17663
rect 23247 17660 23259 17663
rect 23382 17660 23388 17672
rect 23247 17632 23388 17660
rect 23247 17629 23259 17632
rect 23201 17623 23259 17629
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 19978 17552 19984 17604
rect 20036 17592 20042 17604
rect 20625 17595 20683 17601
rect 20625 17592 20637 17595
rect 20036 17564 20637 17592
rect 20036 17552 20042 17564
rect 20625 17561 20637 17564
rect 20671 17561 20683 17595
rect 20625 17555 20683 17561
rect 20714 17552 20720 17604
rect 20772 17592 20778 17604
rect 20809 17595 20867 17601
rect 20809 17592 20821 17595
rect 20772 17564 20821 17592
rect 20772 17552 20778 17564
rect 20809 17561 20821 17564
rect 20855 17561 20867 17595
rect 20809 17555 20867 17561
rect 20993 17595 21051 17601
rect 20993 17561 21005 17595
rect 21039 17592 21051 17595
rect 21269 17595 21327 17601
rect 21269 17592 21281 17595
rect 21039 17564 21281 17592
rect 21039 17561 21051 17564
rect 20993 17555 21051 17561
rect 21269 17561 21281 17564
rect 21315 17561 21327 17595
rect 21269 17555 21327 17561
rect 21358 17552 21364 17604
rect 21416 17552 21422 17604
rect 18414 17524 18420 17536
rect 14884 17496 18420 17524
rect 14884 17484 14890 17496
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 19889 17527 19947 17533
rect 19889 17524 19901 17527
rect 19760 17496 19901 17524
rect 19760 17484 19766 17496
rect 19889 17493 19901 17496
rect 19935 17524 19947 17527
rect 20070 17524 20076 17536
rect 19935 17496 20076 17524
rect 19935 17493 19947 17496
rect 19889 17487 19947 17493
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 21637 17527 21695 17533
rect 21637 17493 21649 17527
rect 21683 17524 21695 17527
rect 22278 17524 22284 17536
rect 21683 17496 22284 17524
rect 21683 17493 21695 17496
rect 21637 17487 21695 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 22738 17484 22744 17536
rect 22796 17484 22802 17536
rect 1104 17434 26312 17456
rect 1104 17382 4761 17434
rect 4813 17382 4825 17434
rect 4877 17382 4889 17434
rect 4941 17382 4953 17434
rect 5005 17382 5017 17434
rect 5069 17382 11063 17434
rect 11115 17382 11127 17434
rect 11179 17382 11191 17434
rect 11243 17382 11255 17434
rect 11307 17382 11319 17434
rect 11371 17382 17365 17434
rect 17417 17382 17429 17434
rect 17481 17382 17493 17434
rect 17545 17382 17557 17434
rect 17609 17382 17621 17434
rect 17673 17382 23667 17434
rect 23719 17382 23731 17434
rect 23783 17382 23795 17434
rect 23847 17382 23859 17434
rect 23911 17382 23923 17434
rect 23975 17382 26312 17434
rect 1104 17360 26312 17382
rect 2406 17280 2412 17332
rect 2464 17320 2470 17332
rect 2501 17323 2559 17329
rect 2501 17320 2513 17323
rect 2464 17292 2513 17320
rect 2464 17280 2470 17292
rect 2501 17289 2513 17292
rect 2547 17289 2559 17323
rect 7466 17320 7472 17332
rect 2501 17283 2559 17289
rect 2746 17292 7472 17320
rect 2225 17255 2283 17261
rect 2225 17221 2237 17255
rect 2271 17252 2283 17255
rect 2746 17252 2774 17292
rect 7466 17280 7472 17292
rect 7524 17280 7530 17332
rect 7576 17292 9168 17320
rect 6178 17252 6184 17264
rect 2271 17224 2774 17252
rect 5934 17224 6184 17252
rect 2271 17221 2283 17224
rect 2225 17215 2283 17221
rect 6178 17212 6184 17224
rect 6236 17212 6242 17264
rect 6365 17255 6423 17261
rect 6365 17221 6377 17255
rect 6411 17221 6423 17255
rect 6365 17215 6423 17221
rect 2130 17144 2136 17196
rect 2188 17144 2194 17196
rect 2314 17144 2320 17196
rect 2372 17184 2378 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 2372 17156 2421 17184
rect 2372 17144 2378 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 4430 17144 4436 17196
rect 4488 17144 4494 17196
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 6052 17182 6224 17184
rect 6385 17182 6413 17215
rect 6454 17212 6460 17264
rect 6512 17252 6518 17264
rect 6565 17255 6623 17261
rect 6565 17252 6577 17255
rect 6512 17224 6577 17252
rect 6512 17212 6518 17224
rect 6565 17221 6577 17224
rect 6611 17221 6623 17255
rect 7576 17252 7604 17292
rect 6565 17215 6623 17221
rect 6748 17224 7604 17252
rect 9140 17252 9168 17292
rect 9306 17280 9312 17332
rect 9364 17280 9370 17332
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 10192 17292 10425 17320
rect 10192 17280 10198 17292
rect 10413 17289 10425 17292
rect 10459 17289 10471 17323
rect 10413 17283 10471 17289
rect 11514 17280 11520 17332
rect 11572 17280 11578 17332
rect 14734 17320 14740 17332
rect 12406 17292 14740 17320
rect 9140 17224 9674 17252
rect 6748 17184 6776 17224
rect 6052 17156 6413 17182
rect 6052 17144 6058 17156
rect 6196 17154 6413 17156
rect 6472 17156 6776 17184
rect 4706 17076 4712 17128
rect 4764 17076 4770 17128
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 5718 17008 5724 17060
rect 5776 17048 5782 17060
rect 6196 17048 6224 17079
rect 6472 17048 6500 17156
rect 6822 17144 6828 17196
rect 6880 17144 6886 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 6932 17156 7573 17184
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 6932 17116 6960 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 8938 17144 8944 17196
rect 8996 17144 9002 17196
rect 9646 17184 9674 17224
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 9824 17224 11008 17252
rect 9824 17212 9830 17224
rect 9646 17156 9996 17184
rect 6604 17088 6960 17116
rect 6604 17076 6610 17088
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7101 17119 7159 17125
rect 7101 17116 7113 17119
rect 7064 17088 7113 17116
rect 7064 17076 7070 17088
rect 7101 17085 7113 17088
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 7837 17119 7895 17125
rect 7837 17085 7849 17119
rect 7883 17116 7895 17119
rect 9030 17116 9036 17128
rect 7883 17088 9036 17116
rect 7883 17085 7895 17088
rect 7837 17079 7895 17085
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 9306 17076 9312 17128
rect 9364 17116 9370 17128
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9364 17088 9873 17116
rect 9364 17076 9370 17088
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 9968 17116 9996 17156
rect 10318 17144 10324 17196
rect 10376 17184 10382 17196
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10376 17156 10609 17184
rect 10376 17144 10382 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10689 17187 10747 17193
rect 10689 17153 10701 17187
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 9968 17088 10456 17116
rect 9861 17079 9919 17085
rect 5776 17020 6500 17048
rect 5776 17008 5782 17020
rect 9950 17008 9956 17060
rect 10008 17048 10014 17060
rect 10137 17051 10195 17057
rect 10137 17048 10149 17051
rect 10008 17020 10149 17048
rect 10008 17008 10014 17020
rect 10137 17017 10149 17020
rect 10183 17017 10195 17051
rect 10137 17011 10195 17017
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 6362 16980 6368 16992
rect 5408 16952 6368 16980
rect 5408 16940 5414 16952
rect 6362 16940 6368 16952
rect 6420 16980 6426 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6420 16952 6561 16980
rect 6420 16940 6426 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 6730 16940 6736 16992
rect 6788 16940 6794 16992
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 6917 16983 6975 16989
rect 6917 16980 6929 16983
rect 6880 16952 6929 16980
rect 6880 16940 6886 16952
rect 6917 16949 6929 16952
rect 6963 16949 6975 16983
rect 6917 16943 6975 16949
rect 7377 16983 7435 16989
rect 7377 16949 7389 16983
rect 7423 16980 7435 16983
rect 8938 16980 8944 16992
rect 7423 16952 8944 16980
rect 7423 16949 7435 16952
rect 7377 16943 7435 16949
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 10284 16952 10333 16980
rect 10284 16940 10290 16952
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 10428 16980 10456 17088
rect 10704 17048 10732 17147
rect 10870 17144 10876 17196
rect 10928 17144 10934 17196
rect 10980 17193 11008 17224
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11664 17156 11713 17184
rect 11664 17144 11670 17156
rect 11701 17153 11713 17156
rect 11747 17184 11759 17187
rect 12406 17184 12434 17292
rect 14734 17280 14740 17292
rect 14792 17280 14798 17332
rect 18230 17320 18236 17332
rect 16316 17292 18236 17320
rect 13909 17255 13967 17261
rect 13909 17221 13921 17255
rect 13955 17221 13967 17255
rect 13909 17215 13967 17221
rect 11747 17156 12434 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 11790 17076 11796 17128
rect 11848 17076 11854 17128
rect 11882 17076 11888 17128
rect 11940 17076 11946 17128
rect 11977 17119 12035 17125
rect 11977 17085 11989 17119
rect 12023 17116 12035 17119
rect 12710 17116 12716 17128
rect 12023 17088 12716 17116
rect 12023 17085 12035 17088
rect 11977 17079 12035 17085
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 13924 17116 13952 17215
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 14109 17255 14167 17261
rect 14109 17252 14121 17255
rect 14056 17224 14121 17252
rect 14056 17212 14062 17224
rect 14109 17221 14121 17224
rect 14155 17221 14167 17255
rect 14109 17215 14167 17221
rect 14550 17144 14556 17196
rect 14608 17144 14614 17196
rect 16316 17193 16344 17292
rect 18230 17280 18236 17292
rect 18288 17280 18294 17332
rect 18414 17280 18420 17332
rect 18472 17280 18478 17332
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 21545 17323 21603 17329
rect 21545 17320 21557 17323
rect 21324 17292 21557 17320
rect 21324 17280 21330 17292
rect 21545 17289 21557 17292
rect 21591 17289 21603 17323
rect 21545 17283 21603 17289
rect 21652 17292 24072 17320
rect 16393 17255 16451 17261
rect 16393 17221 16405 17255
rect 16439 17252 16451 17255
rect 16945 17255 17003 17261
rect 16945 17252 16957 17255
rect 16439 17224 16957 17252
rect 16439 17221 16451 17224
rect 16393 17215 16451 17221
rect 16945 17221 16957 17224
rect 16991 17221 17003 17255
rect 16945 17215 17003 17221
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 21652 17252 21680 17292
rect 20456 17224 21680 17252
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17184 19671 17187
rect 19794 17184 19800 17196
rect 19659 17156 19800 17184
rect 19659 17153 19671 17156
rect 19613 17147 19671 17153
rect 14182 17116 14188 17128
rect 13924 17088 14188 17116
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 14844 17116 14872 17147
rect 19794 17144 19800 17156
rect 19852 17184 19858 17196
rect 20456 17193 20484 17224
rect 22278 17212 22284 17264
rect 22336 17212 22342 17264
rect 24044 17261 24072 17292
rect 24029 17255 24087 17261
rect 24029 17221 24041 17255
rect 24075 17221 24087 17255
rect 24029 17215 24087 17221
rect 20441 17187 20499 17193
rect 20441 17184 20453 17187
rect 19852 17156 20453 17184
rect 19852 17144 19858 17156
rect 20441 17153 20453 17156
rect 20487 17153 20499 17187
rect 21450 17184 21456 17196
rect 20441 17147 20499 17153
rect 20824 17156 21456 17184
rect 14292 17088 14872 17116
rect 13630 17048 13636 17060
rect 10704 17020 13636 17048
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 14292 17057 14320 17088
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 16632 17088 16681 17116
rect 16632 17076 16638 17088
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 14277 17051 14335 17057
rect 14277 17017 14289 17051
rect 14323 17017 14335 17051
rect 19720 17048 19748 17079
rect 19978 17076 19984 17128
rect 20036 17076 20042 17128
rect 20530 17076 20536 17128
rect 20588 17076 20594 17128
rect 20824 17125 20852 17156
rect 21450 17144 21456 17156
rect 21508 17144 21514 17196
rect 22002 17144 22008 17196
rect 22060 17144 22066 17196
rect 23414 17156 23520 17184
rect 23492 17128 23520 17156
rect 25682 17144 25688 17196
rect 25740 17144 25746 17196
rect 20809 17119 20867 17125
rect 20809 17085 20821 17119
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 20990 17076 20996 17128
rect 21048 17076 21054 17128
rect 23474 17076 23480 17128
rect 23532 17076 23538 17128
rect 20070 17048 20076 17060
rect 19720 17020 20076 17048
rect 14277 17011 14335 17017
rect 20070 17008 20076 17020
rect 20128 17008 20134 17060
rect 25866 17008 25872 17060
rect 25924 17008 25930 17060
rect 10870 16980 10876 16992
rect 10428 16952 10876 16980
rect 10321 16943 10379 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16980 14151 16983
rect 14182 16980 14188 16992
rect 14139 16952 14188 16980
rect 14139 16949 14151 16952
rect 14093 16943 14151 16949
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 14737 16983 14795 16989
rect 14737 16980 14749 16983
rect 14700 16952 14749 16980
rect 14700 16940 14706 16952
rect 14737 16949 14749 16952
rect 14783 16949 14795 16983
rect 14737 16943 14795 16949
rect 15013 16983 15071 16989
rect 15013 16949 15025 16983
rect 15059 16980 15071 16983
rect 15102 16980 15108 16992
rect 15059 16952 15108 16980
rect 15059 16949 15071 16952
rect 15013 16943 15071 16949
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 20898 16980 20904 16992
rect 18564 16952 20904 16980
rect 18564 16940 18570 16952
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 1104 16890 26312 16912
rect 1104 16838 4101 16890
rect 4153 16838 4165 16890
rect 4217 16838 4229 16890
rect 4281 16838 4293 16890
rect 4345 16838 4357 16890
rect 4409 16838 10403 16890
rect 10455 16838 10467 16890
rect 10519 16838 10531 16890
rect 10583 16838 10595 16890
rect 10647 16838 10659 16890
rect 10711 16838 16705 16890
rect 16757 16838 16769 16890
rect 16821 16838 16833 16890
rect 16885 16838 16897 16890
rect 16949 16838 16961 16890
rect 17013 16838 23007 16890
rect 23059 16838 23071 16890
rect 23123 16838 23135 16890
rect 23187 16838 23199 16890
rect 23251 16838 23263 16890
rect 23315 16838 26312 16890
rect 1104 16816 26312 16838
rect 1397 16779 1455 16785
rect 1397 16745 1409 16779
rect 1443 16776 1455 16779
rect 2130 16776 2136 16788
rect 1443 16748 2136 16776
rect 1443 16745 1455 16748
rect 1397 16739 1455 16745
rect 2130 16736 2136 16748
rect 2188 16736 2194 16788
rect 4614 16736 4620 16788
rect 4672 16736 4678 16788
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 4985 16779 5043 16785
rect 4985 16776 4997 16779
rect 4764 16748 4997 16776
rect 4764 16736 4770 16748
rect 4985 16745 4997 16748
rect 5031 16745 5043 16779
rect 4985 16739 5043 16745
rect 6086 16736 6092 16788
rect 6144 16776 6150 16788
rect 6822 16776 6828 16788
rect 6144 16748 6828 16776
rect 6144 16736 6150 16748
rect 6822 16736 6828 16748
rect 6880 16776 6886 16788
rect 6880 16748 7144 16776
rect 6880 16736 6886 16748
rect 6454 16708 6460 16720
rect 4356 16680 6460 16708
rect 934 16532 940 16584
rect 992 16572 998 16584
rect 4356 16581 4384 16680
rect 6454 16668 6460 16680
rect 6512 16668 6518 16720
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16640 4675 16643
rect 5810 16640 5816 16652
rect 4663 16612 5816 16640
rect 4663 16609 4675 16612
rect 4617 16603 4675 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6270 16640 6276 16652
rect 5951 16612 6276 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 6604 16612 7021 16640
rect 6604 16600 6610 16612
rect 7009 16609 7021 16612
rect 7055 16609 7067 16643
rect 7116 16640 7144 16748
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 8720 16748 8769 16776
rect 8720 16736 8726 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 13909 16779 13967 16785
rect 8757 16739 8815 16745
rect 11992 16748 12296 16776
rect 8772 16640 8800 16739
rect 9122 16668 9128 16720
rect 9180 16708 9186 16720
rect 9950 16708 9956 16720
rect 9180 16680 9956 16708
rect 9180 16668 9186 16680
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 10042 16668 10048 16720
rect 10100 16708 10106 16720
rect 10689 16711 10747 16717
rect 10100 16680 10640 16708
rect 10100 16668 10106 16680
rect 7116 16612 8708 16640
rect 8772 16612 9812 16640
rect 7009 16603 7067 16609
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 992 16544 1593 16572
rect 992 16532 998 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 1581 16535 1639 16541
rect 4341 16575 4399 16581
rect 4341 16541 4353 16575
rect 4387 16541 4399 16575
rect 4341 16535 4399 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16572 5227 16575
rect 5629 16575 5687 16581
rect 5215 16544 5304 16572
rect 5215 16541 5227 16544
rect 5169 16535 5227 16541
rect 3970 16396 3976 16448
rect 4028 16436 4034 16448
rect 5276 16445 5304 16544
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 5718 16572 5724 16584
rect 5675 16544 5724 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 5718 16532 5724 16544
rect 5776 16532 5782 16584
rect 6086 16532 6092 16584
rect 6144 16532 6150 16584
rect 6178 16532 6184 16584
rect 6236 16532 6242 16584
rect 8680 16572 8708 16612
rect 9784 16584 9812 16612
rect 10318 16600 10324 16652
rect 10376 16600 10382 16652
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 8680 16544 8953 16572
rect 8941 16541 8953 16544
rect 8987 16572 8999 16575
rect 9122 16572 9128 16584
rect 8987 16544 9128 16572
rect 8987 16541 8999 16544
rect 8941 16535 8999 16541
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9766 16532 9772 16584
rect 9824 16532 9830 16584
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 10045 16575 10103 16581
rect 10045 16572 10057 16575
rect 9907 16544 10057 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 10045 16541 10057 16544
rect 10091 16541 10103 16575
rect 10045 16535 10103 16541
rect 10193 16575 10251 16581
rect 10193 16541 10205 16575
rect 10239 16572 10251 16575
rect 10336 16572 10364 16600
rect 10510 16575 10568 16581
rect 10510 16572 10522 16575
rect 10239 16541 10272 16572
rect 10336 16544 10522 16572
rect 10193 16535 10272 16541
rect 10510 16541 10522 16544
rect 10556 16541 10568 16575
rect 10510 16535 10568 16541
rect 7282 16464 7288 16516
rect 7340 16464 7346 16516
rect 9033 16507 9091 16513
rect 9033 16504 9045 16507
rect 8510 16476 9045 16504
rect 9033 16473 9045 16476
rect 9079 16473 9091 16507
rect 9033 16467 9091 16473
rect 4893 16439 4951 16445
rect 4893 16436 4905 16439
rect 4028 16408 4905 16436
rect 4028 16396 4034 16408
rect 4893 16405 4905 16408
rect 4939 16405 4951 16439
rect 4893 16399 4951 16405
rect 5261 16439 5319 16445
rect 5261 16405 5273 16439
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 5721 16439 5779 16445
rect 5721 16436 5733 16439
rect 5592 16408 5733 16436
rect 5592 16396 5598 16408
rect 5721 16405 5733 16408
rect 5767 16436 5779 16439
rect 6638 16436 6644 16448
rect 5767 16408 6644 16436
rect 5767 16405 5779 16408
rect 5721 16399 5779 16405
rect 6638 16396 6644 16408
rect 6696 16396 6702 16448
rect 10244 16436 10272 16535
rect 10318 16464 10324 16516
rect 10376 16464 10382 16516
rect 10413 16507 10471 16513
rect 10413 16473 10425 16507
rect 10459 16504 10471 16507
rect 10612 16504 10640 16680
rect 10689 16677 10701 16711
rect 10735 16708 10747 16711
rect 10735 16680 11928 16708
rect 10735 16677 10747 16680
rect 10689 16671 10747 16677
rect 11149 16643 11207 16649
rect 11149 16609 11161 16643
rect 11195 16640 11207 16643
rect 11330 16640 11336 16652
rect 11195 16612 11336 16640
rect 11195 16609 11207 16612
rect 11149 16603 11207 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11422 16600 11428 16652
rect 11480 16600 11486 16652
rect 11514 16532 11520 16584
rect 11572 16532 11578 16584
rect 11900 16581 11928 16680
rect 11992 16640 12020 16748
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 12124 16680 12204 16708
rect 12124 16668 12130 16680
rect 12176 16649 12204 16680
rect 12161 16643 12219 16649
rect 11992 16612 12112 16640
rect 12084 16581 12112 16612
rect 12161 16609 12173 16643
rect 12207 16609 12219 16643
rect 12268 16640 12296 16748
rect 13909 16745 13921 16779
rect 13955 16776 13967 16779
rect 13998 16776 14004 16788
rect 13955 16748 14004 16776
rect 13955 16745 13967 16748
rect 13909 16739 13967 16745
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 20714 16776 20720 16788
rect 19720 16748 20720 16776
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 18506 16708 18512 16720
rect 13688 16680 18512 16708
rect 13688 16668 13694 16680
rect 18506 16668 18512 16680
rect 18564 16668 18570 16720
rect 13446 16640 13452 16652
rect 12268 16612 13452 16640
rect 12161 16603 12219 16609
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 14366 16640 14372 16652
rect 14108 16612 14372 16640
rect 14108 16581 14136 16612
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 19720 16640 19748 16748
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 20898 16736 20904 16788
rect 20956 16776 20962 16788
rect 25682 16776 25688 16788
rect 20956 16748 25688 16776
rect 20956 16736 20962 16748
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 19797 16711 19855 16717
rect 19797 16677 19809 16711
rect 19843 16708 19855 16711
rect 20806 16708 20812 16720
rect 19843 16680 20812 16708
rect 19843 16677 19855 16680
rect 19797 16671 19855 16677
rect 20806 16668 20812 16680
rect 20864 16668 20870 16720
rect 23198 16668 23204 16720
rect 23256 16668 23262 16720
rect 19720 16612 19840 16640
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16541 11943 16575
rect 11885 16535 11943 16541
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 17221 16575 17279 16581
rect 17221 16572 17233 16575
rect 15620 16544 17233 16572
rect 15620 16532 15626 16544
rect 17221 16541 17233 16544
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 17313 16575 17371 16581
rect 17313 16541 17325 16575
rect 17359 16572 17371 16575
rect 17954 16572 17960 16584
rect 17359 16544 17960 16572
rect 17359 16541 17371 16544
rect 17313 16535 17371 16541
rect 10459 16476 10640 16504
rect 10459 16473 10471 16476
rect 10413 16467 10471 16473
rect 12434 16464 12440 16516
rect 12492 16464 12498 16516
rect 14185 16507 14243 16513
rect 14185 16504 14197 16507
rect 13662 16476 14197 16504
rect 14185 16473 14197 16476
rect 14231 16473 14243 16507
rect 17236 16504 17264 16535
rect 17954 16532 17960 16544
rect 18012 16532 18018 16584
rect 19812 16581 19840 16612
rect 19886 16600 19892 16652
rect 19944 16640 19950 16652
rect 20165 16643 20223 16649
rect 19944 16612 20116 16640
rect 19944 16600 19950 16612
rect 20088 16581 20116 16612
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 21358 16640 21364 16652
rect 20211 16612 20576 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 20548 16584 20576 16612
rect 21106 16612 21364 16640
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16541 20131 16575
rect 20073 16535 20131 16541
rect 18046 16504 18052 16516
rect 17236 16476 18052 16504
rect 14185 16467 14243 16473
rect 18046 16464 18052 16476
rect 18104 16464 18110 16516
rect 12066 16436 12072 16448
rect 10244 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 19996 16436 20024 16535
rect 20254 16532 20260 16584
rect 20312 16532 20318 16584
rect 20530 16532 20536 16584
rect 20588 16532 20594 16584
rect 20714 16532 20720 16584
rect 20772 16532 20778 16584
rect 21106 16574 21134 16612
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 21450 16600 21456 16652
rect 21508 16640 21514 16652
rect 22094 16640 22100 16652
rect 21508 16612 22100 16640
rect 21508 16600 21514 16612
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 23566 16640 23572 16652
rect 23400 16612 23572 16640
rect 21177 16575 21235 16581
rect 21177 16574 21189 16575
rect 21106 16572 21189 16574
rect 20916 16546 21189 16572
rect 20916 16544 21134 16546
rect 20162 16464 20168 16516
rect 20220 16504 20226 16516
rect 20349 16507 20407 16513
rect 20349 16504 20361 16507
rect 20220 16476 20361 16504
rect 20220 16464 20226 16476
rect 20349 16473 20361 16476
rect 20395 16473 20407 16507
rect 20349 16467 20407 16473
rect 20916 16436 20944 16544
rect 21177 16541 21189 16546
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 21266 16532 21272 16584
rect 21324 16532 21330 16584
rect 23400 16581 23428 16612
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16574 23443 16575
rect 23431 16546 23465 16574
rect 23431 16541 23443 16546
rect 23385 16535 23443 16541
rect 20990 16464 20996 16516
rect 21048 16464 21054 16516
rect 21729 16507 21787 16513
rect 21729 16473 21741 16507
rect 21775 16504 21787 16507
rect 21818 16504 21824 16516
rect 21775 16476 21824 16504
rect 21775 16473 21787 16476
rect 21729 16467 21787 16473
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 22738 16464 22744 16516
rect 22796 16464 22802 16516
rect 19996 16408 20944 16436
rect 21082 16396 21088 16448
rect 21140 16445 21146 16448
rect 21140 16399 21149 16445
rect 21140 16396 21146 16399
rect 23474 16396 23480 16448
rect 23532 16396 23538 16448
rect 1104 16346 26312 16368
rect 1104 16294 4761 16346
rect 4813 16294 4825 16346
rect 4877 16294 4889 16346
rect 4941 16294 4953 16346
rect 5005 16294 5017 16346
rect 5069 16294 11063 16346
rect 11115 16294 11127 16346
rect 11179 16294 11191 16346
rect 11243 16294 11255 16346
rect 11307 16294 11319 16346
rect 11371 16294 17365 16346
rect 17417 16294 17429 16346
rect 17481 16294 17493 16346
rect 17545 16294 17557 16346
rect 17609 16294 17621 16346
rect 17673 16294 23667 16346
rect 23719 16294 23731 16346
rect 23783 16294 23795 16346
rect 23847 16294 23859 16346
rect 23911 16294 23923 16346
rect 23975 16294 26312 16346
rect 1104 16272 26312 16294
rect 2314 16192 2320 16244
rect 2372 16192 2378 16244
rect 3329 16235 3387 16241
rect 3329 16201 3341 16235
rect 3375 16201 3387 16235
rect 3329 16195 3387 16201
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3786 16232 3792 16244
rect 3743 16204 3792 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 2332 16164 2360 16192
rect 3344 16164 3372 16195
rect 3786 16192 3792 16204
rect 3844 16232 3850 16244
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 3844 16204 5365 16232
rect 3844 16192 3850 16204
rect 5353 16201 5365 16204
rect 5399 16232 5411 16235
rect 5399 16204 6132 16232
rect 5399 16201 5411 16204
rect 5353 16195 5411 16201
rect 2332 16136 2774 16164
rect 2314 16056 2320 16108
rect 2372 16056 2378 16108
rect 2424 16105 2452 16136
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16065 2467 16099
rect 2409 16059 2467 16065
rect 2746 16028 2774 16136
rect 2884 16136 3372 16164
rect 2884 16105 2912 16136
rect 5442 16124 5448 16176
rect 5500 16124 5506 16176
rect 6104 16164 6132 16204
rect 6638 16192 6644 16244
rect 6696 16232 6702 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6696 16204 6837 16232
rect 6696 16192 6702 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 6825 16195 6883 16201
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7340 16204 8217 16232
rect 7340 16192 7346 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 10318 16192 10324 16244
rect 10376 16192 10382 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16232 10563 16235
rect 11514 16232 11520 16244
rect 10551 16204 11520 16232
rect 10551 16201 10563 16204
rect 10505 16195 10563 16201
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 12710 16192 12716 16244
rect 12768 16192 12774 16244
rect 13446 16192 13452 16244
rect 13504 16192 13510 16244
rect 19242 16232 19248 16244
rect 16960 16204 19248 16232
rect 8570 16164 8576 16176
rect 6104 16136 8576 16164
rect 8570 16124 8576 16136
rect 8628 16124 8634 16176
rect 10336 16164 10364 16192
rect 12345 16167 12403 16173
rect 12345 16164 12357 16167
rect 10336 16136 12357 16164
rect 12345 16133 12357 16136
rect 12391 16133 12403 16167
rect 12345 16127 12403 16133
rect 12437 16167 12495 16173
rect 12437 16133 12449 16167
rect 12483 16164 12495 16167
rect 15102 16164 15108 16176
rect 12483 16136 15108 16164
rect 12483 16133 12495 16136
rect 12437 16127 12495 16133
rect 15102 16124 15108 16136
rect 15160 16124 15166 16176
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16096 3019 16099
rect 5460 16096 5488 16124
rect 6733 16099 6791 16105
rect 3007 16068 4108 16096
rect 5460 16068 5580 16096
rect 3007 16065 3019 16068
rect 2961 16059 3019 16065
rect 2976 16028 3004 16059
rect 2746 16000 3004 16028
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 16028 3847 16031
rect 3878 16028 3884 16040
rect 3835 16000 3884 16028
rect 3835 15997 3847 16000
rect 3789 15991 3847 15997
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 3970 15988 3976 16040
rect 4028 15988 4034 16040
rect 2501 15963 2559 15969
rect 2501 15929 2513 15963
rect 2547 15960 2559 15963
rect 2774 15960 2780 15972
rect 2547 15932 2780 15960
rect 2547 15929 2559 15932
rect 2501 15923 2559 15929
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 4080 15960 4108 16068
rect 5442 15988 5448 16040
rect 5500 15988 5506 16040
rect 5552 16037 5580 16068
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 6779 16068 8125 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 8113 16065 8125 16068
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 8386 16056 8392 16108
rect 8444 16056 8450 16108
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10229 16099 10287 16105
rect 10229 16096 10241 16099
rect 9824 16068 10241 16096
rect 9824 16056 9830 16068
rect 10229 16065 10241 16068
rect 10275 16065 10287 16099
rect 10229 16059 10287 16065
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 10778 16096 10784 16108
rect 10367 16068 10784 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 15997 5595 16031
rect 5537 15991 5595 15997
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 4080 15932 5304 15960
rect 1670 15852 1676 15904
rect 1728 15892 1734 15904
rect 2133 15895 2191 15901
rect 2133 15892 2145 15895
rect 1728 15864 2145 15892
rect 1728 15852 1734 15864
rect 2133 15861 2145 15864
rect 2179 15861 2191 15895
rect 2133 15855 2191 15861
rect 2222 15852 2228 15904
rect 2280 15892 2286 15904
rect 2685 15895 2743 15901
rect 2685 15892 2697 15895
rect 2280 15864 2697 15892
rect 2280 15852 2286 15864
rect 2685 15861 2697 15864
rect 2731 15861 2743 15895
rect 2685 15855 2743 15861
rect 2958 15852 2964 15904
rect 3016 15892 3022 15904
rect 3053 15895 3111 15901
rect 3053 15892 3065 15895
rect 3016 15864 3065 15892
rect 3016 15852 3022 15864
rect 3053 15861 3065 15864
rect 3099 15861 3111 15895
rect 3053 15855 3111 15861
rect 4985 15895 5043 15901
rect 4985 15861 4997 15895
rect 5031 15892 5043 15895
rect 5166 15892 5172 15904
rect 5031 15864 5172 15892
rect 5031 15861 5043 15864
rect 4985 15855 5043 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5276 15892 5304 15932
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 6932 15960 6960 15991
rect 7558 15988 7564 16040
rect 7616 15988 7622 16040
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 10870 16028 10876 16040
rect 10551 16000 10876 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 12176 16028 12204 16059
rect 12526 16056 12532 16108
rect 12584 16096 12590 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 12584 16068 13277 16096
rect 12584 16056 12590 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16960 16105 16988 16204
rect 19242 16192 19248 16204
rect 19300 16232 19306 16244
rect 20349 16235 20407 16241
rect 20349 16232 20361 16235
rect 19300 16204 20361 16232
rect 19300 16192 19306 16204
rect 20349 16201 20361 16204
rect 20395 16232 20407 16235
rect 20714 16232 20720 16244
rect 20395 16204 20720 16232
rect 20395 16201 20407 16204
rect 20349 16195 20407 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 21545 16235 21603 16241
rect 21545 16232 21557 16235
rect 21232 16204 21557 16232
rect 21232 16192 21238 16204
rect 21545 16201 21557 16204
rect 21591 16201 21603 16235
rect 21545 16195 21603 16201
rect 18230 16124 18236 16176
rect 18288 16124 18294 16176
rect 19058 16124 19064 16176
rect 19116 16124 19122 16176
rect 21082 16124 21088 16176
rect 21140 16164 21146 16176
rect 21821 16167 21879 16173
rect 21821 16164 21833 16167
rect 21140 16136 21833 16164
rect 21140 16124 21146 16136
rect 21821 16133 21833 16136
rect 21867 16133 21879 16167
rect 21821 16127 21879 16133
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16632 16068 16957 16096
rect 16632 16056 16638 16068
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 20864 16068 22017 16096
rect 20864 16056 20870 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22097 16099 22155 16105
rect 22097 16065 22109 16099
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 12710 16028 12716 16040
rect 12176 16000 12716 16028
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 16028 13139 16031
rect 14642 16028 14648 16040
rect 13127 16000 14648 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17770 16028 17776 16040
rect 17267 16000 17776 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 6788 15932 6960 15960
rect 6788 15920 6794 15932
rect 5994 15892 6000 15904
rect 5276 15864 6000 15892
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6362 15852 6368 15904
rect 6420 15852 6426 15904
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 18984 15892 19012 15991
rect 20990 15988 20996 16040
rect 21048 15988 21054 16040
rect 21266 15988 21272 16040
rect 21324 16028 21330 16040
rect 22112 16028 22140 16059
rect 21324 16000 22140 16028
rect 21324 15988 21330 16000
rect 21818 15920 21824 15972
rect 21876 15920 21882 15972
rect 17092 15864 19012 15892
rect 17092 15852 17098 15864
rect 1104 15802 26312 15824
rect 1104 15750 4101 15802
rect 4153 15750 4165 15802
rect 4217 15750 4229 15802
rect 4281 15750 4293 15802
rect 4345 15750 4357 15802
rect 4409 15750 10403 15802
rect 10455 15750 10467 15802
rect 10519 15750 10531 15802
rect 10583 15750 10595 15802
rect 10647 15750 10659 15802
rect 10711 15750 16705 15802
rect 16757 15750 16769 15802
rect 16821 15750 16833 15802
rect 16885 15750 16897 15802
rect 16949 15750 16961 15802
rect 17013 15750 23007 15802
rect 23059 15750 23071 15802
rect 23123 15750 23135 15802
rect 23187 15750 23199 15802
rect 23251 15750 23263 15802
rect 23315 15750 26312 15802
rect 1104 15728 26312 15750
rect 2314 15648 2320 15700
rect 2372 15688 2378 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 2372 15660 3801 15688
rect 2372 15648 2378 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 5994 15648 6000 15700
rect 6052 15688 6058 15700
rect 7926 15688 7932 15700
rect 6052 15660 7932 15688
rect 6052 15648 6058 15660
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 11885 15691 11943 15697
rect 11885 15657 11897 15691
rect 11931 15688 11943 15691
rect 12434 15688 12440 15700
rect 11931 15660 12440 15688
rect 11931 15657 11943 15660
rect 11885 15651 11943 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 16485 15691 16543 15697
rect 16485 15657 16497 15691
rect 16531 15688 16543 15691
rect 17586 15688 17592 15700
rect 16531 15660 17592 15688
rect 16531 15657 16543 15660
rect 16485 15651 16543 15657
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 17770 15648 17776 15700
rect 17828 15648 17834 15700
rect 18141 15691 18199 15697
rect 18141 15657 18153 15691
rect 18187 15688 18199 15691
rect 18230 15688 18236 15700
rect 18187 15660 18236 15688
rect 18187 15657 18199 15660
rect 18141 15651 18199 15657
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 20990 15648 20996 15700
rect 21048 15688 21054 15700
rect 22143 15691 22201 15697
rect 22143 15688 22155 15691
rect 21048 15660 22155 15688
rect 21048 15648 21054 15660
rect 22143 15657 22155 15660
rect 22189 15657 22201 15691
rect 22143 15651 22201 15657
rect 3329 15623 3387 15629
rect 3329 15589 3341 15623
rect 3375 15620 3387 15623
rect 3878 15620 3884 15632
rect 3375 15592 3884 15620
rect 3375 15589 3387 15592
rect 3329 15583 3387 15589
rect 3878 15580 3884 15592
rect 3936 15620 3942 15632
rect 6454 15620 6460 15632
rect 3936 15592 6460 15620
rect 3936 15580 3942 15592
rect 6454 15580 6460 15592
rect 6512 15580 6518 15632
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 19058 15620 19064 15632
rect 13780 15592 19064 15620
rect 13780 15580 13786 15592
rect 19058 15580 19064 15592
rect 19116 15580 19122 15632
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 1581 15555 1639 15561
rect 1581 15552 1593 15555
rect 1452 15524 1593 15552
rect 1452 15512 1458 15524
rect 1581 15521 1593 15524
rect 1627 15521 1639 15555
rect 1581 15515 1639 15521
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 2222 15552 2228 15564
rect 1903 15524 2228 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4522 15552 4528 15564
rect 4479 15524 4528 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 7374 15512 7380 15564
rect 7432 15552 7438 15564
rect 7653 15555 7711 15561
rect 7653 15552 7665 15555
rect 7432 15524 7665 15552
rect 7432 15512 7438 15524
rect 7653 15521 7665 15524
rect 7699 15521 7711 15555
rect 15470 15552 15476 15564
rect 7653 15515 7711 15521
rect 7852 15524 15476 15552
rect 2958 15444 2964 15496
rect 3016 15444 3022 15496
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 3844 15456 4169 15484
rect 3844 15444 3850 15456
rect 4157 15453 4169 15456
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 5258 15444 5264 15496
rect 5316 15444 5322 15496
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15484 7619 15487
rect 7852 15484 7880 15524
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 15930 15512 15936 15564
rect 15988 15552 15994 15564
rect 16025 15555 16083 15561
rect 16025 15552 16037 15555
rect 15988 15524 16037 15552
rect 15988 15512 15994 15524
rect 16025 15521 16037 15524
rect 16071 15521 16083 15555
rect 16025 15515 16083 15521
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 16942 15552 16948 15564
rect 16899 15524 16948 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 17034 15512 17040 15564
rect 17092 15512 17098 15564
rect 17126 15512 17132 15564
rect 17184 15512 17190 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 18064 15524 19441 15552
rect 7607 15456 7880 15484
rect 7607 15453 7619 15456
rect 7561 15447 7619 15453
rect 7926 15444 7932 15496
rect 7984 15444 7990 15496
rect 8110 15444 8116 15496
rect 8168 15484 8174 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8168 15456 8953 15484
rect 8168 15444 8174 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 10008 15456 10057 15484
rect 10008 15444 10014 15456
rect 10045 15453 10057 15456
rect 10091 15484 10103 15487
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 10091 15456 10333 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10321 15453 10333 15456
rect 10367 15453 10379 15487
rect 10321 15447 10379 15453
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12069 15487 12127 15493
rect 12069 15484 12081 15487
rect 11940 15456 12081 15484
rect 11940 15444 11946 15456
rect 12069 15453 12081 15456
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 14458 15484 14464 15496
rect 13587 15456 14464 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 15562 15444 15568 15496
rect 15620 15444 15626 15496
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15484 16175 15487
rect 16482 15484 16488 15496
rect 16163 15456 16488 15484
rect 16163 15453 16175 15456
rect 16117 15447 16175 15453
rect 16482 15444 16488 15456
rect 16540 15484 16546 15496
rect 16761 15487 16819 15493
rect 16761 15484 16773 15487
rect 16540 15456 16773 15484
rect 16540 15444 16546 15456
rect 16761 15453 16773 15456
rect 16807 15484 16819 15487
rect 17052 15484 17080 15512
rect 18064 15496 18092 15524
rect 19429 15521 19441 15524
rect 19475 15552 19487 15555
rect 19978 15552 19984 15564
rect 19475 15524 19984 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 20349 15555 20407 15561
rect 20349 15521 20361 15555
rect 20395 15552 20407 15555
rect 20622 15552 20628 15564
rect 20395 15524 20628 15552
rect 20395 15521 20407 15524
rect 20349 15515 20407 15521
rect 20622 15512 20628 15524
rect 20680 15552 20686 15564
rect 21450 15552 21456 15564
rect 20680 15524 21456 15552
rect 20680 15512 20686 15524
rect 21450 15512 21456 15524
rect 21508 15512 21514 15564
rect 16807 15456 17080 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 17218 15444 17224 15496
rect 17276 15444 17282 15496
rect 17586 15444 17592 15496
rect 17644 15444 17650 15496
rect 18046 15444 18052 15496
rect 18104 15444 18110 15496
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 19208 15456 19257 15484
rect 19208 15444 19214 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 20806 15484 20812 15496
rect 20763 15456 20812 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 7469 15419 7527 15425
rect 7469 15385 7481 15419
rect 7515 15416 7527 15419
rect 8570 15416 8576 15428
rect 7515 15388 8576 15416
rect 7515 15385 7527 15388
rect 7469 15379 7527 15385
rect 8570 15376 8576 15388
rect 8628 15376 8634 15428
rect 17034 15376 17040 15428
rect 17092 15416 17098 15428
rect 17405 15419 17463 15425
rect 17405 15416 17417 15419
rect 17092 15388 17417 15416
rect 17092 15376 17098 15388
rect 17405 15385 17417 15388
rect 17451 15385 17463 15419
rect 17405 15379 17463 15385
rect 17497 15419 17555 15425
rect 17497 15385 17509 15419
rect 17543 15416 17555 15419
rect 17862 15416 17868 15428
rect 17543 15388 17868 15416
rect 17543 15385 17555 15388
rect 17497 15379 17555 15385
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 4249 15351 4307 15357
rect 4249 15317 4261 15351
rect 4295 15348 4307 15351
rect 4522 15348 4528 15360
rect 4295 15320 4528 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 6546 15308 6552 15360
rect 6604 15308 6610 15360
rect 7101 15351 7159 15357
rect 7101 15317 7113 15351
rect 7147 15348 7159 15351
rect 7282 15348 7288 15360
rect 7147 15320 7288 15348
rect 7147 15317 7159 15320
rect 7101 15311 7159 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15348 8079 15351
rect 8294 15348 8300 15360
rect 8067 15320 8300 15348
rect 8067 15317 8079 15320
rect 8021 15311 8079 15317
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 9585 15351 9643 15357
rect 9585 15348 9597 15351
rect 9364 15320 9597 15348
rect 9364 15308 9370 15320
rect 9585 15317 9597 15320
rect 9631 15317 9643 15351
rect 9585 15311 9643 15317
rect 9677 15351 9735 15357
rect 9677 15317 9689 15351
rect 9723 15348 9735 15351
rect 9766 15348 9772 15360
rect 9723 15320 9772 15348
rect 9723 15317 9735 15320
rect 9677 15311 9735 15317
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 10134 15308 10140 15360
rect 10192 15308 10198 15360
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10413 15351 10471 15357
rect 10413 15348 10425 15351
rect 10284 15320 10425 15348
rect 10284 15308 10290 15320
rect 10413 15317 10425 15320
rect 10459 15317 10471 15351
rect 10413 15311 10471 15317
rect 13630 15308 13636 15360
rect 13688 15348 13694 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13688 15320 13737 15348
rect 13688 15308 13694 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 15657 15351 15715 15357
rect 15657 15317 15669 15351
rect 15703 15348 15715 15351
rect 15746 15348 15752 15360
rect 15703 15320 15752 15348
rect 15703 15317 15715 15320
rect 15657 15311 15715 15317
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 17678 15348 17684 15360
rect 16908 15320 17684 15348
rect 16908 15308 16914 15320
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 19260 15348 19288 15447
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 21082 15376 21088 15428
rect 21140 15376 21146 15428
rect 23382 15348 23388 15360
rect 19260 15320 23388 15348
rect 23382 15308 23388 15320
rect 23440 15348 23446 15360
rect 24302 15348 24308 15360
rect 23440 15320 24308 15348
rect 23440 15308 23446 15320
rect 24302 15308 24308 15320
rect 24360 15308 24366 15360
rect 1104 15258 26312 15280
rect 1104 15206 4761 15258
rect 4813 15206 4825 15258
rect 4877 15206 4889 15258
rect 4941 15206 4953 15258
rect 5005 15206 5017 15258
rect 5069 15206 11063 15258
rect 11115 15206 11127 15258
rect 11179 15206 11191 15258
rect 11243 15206 11255 15258
rect 11307 15206 11319 15258
rect 11371 15206 17365 15258
rect 17417 15206 17429 15258
rect 17481 15206 17493 15258
rect 17545 15206 17557 15258
rect 17609 15206 17621 15258
rect 17673 15206 23667 15258
rect 23719 15206 23731 15258
rect 23783 15206 23795 15258
rect 23847 15206 23859 15258
rect 23911 15206 23923 15258
rect 23975 15206 26312 15258
rect 1104 15184 26312 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 6546 15144 6552 15156
rect 1452 15116 6552 15144
rect 1452 15104 1458 15116
rect 1670 15036 1676 15088
rect 1728 15036 1734 15088
rect 1394 14968 1400 15020
rect 1452 14968 1458 15020
rect 2774 14968 2780 15020
rect 2832 14968 2838 15020
rect 4172 15017 4200 15116
rect 5718 15076 5724 15088
rect 5658 15048 5724 15076
rect 5718 15036 5724 15048
rect 5776 15036 5782 15088
rect 6380 15017 6408 15116
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 8110 15144 8116 15156
rect 7616 15116 8116 15144
rect 7616 15104 7622 15116
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8220 15116 10824 15144
rect 7098 15036 7104 15088
rect 7156 15036 7162 15088
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14940 4491 14943
rect 4890 14940 4896 14952
rect 4479 14912 4896 14940
rect 4479 14909 4491 14912
rect 4433 14903 4491 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5442 14900 5448 14952
rect 5500 14940 5506 14952
rect 6181 14943 6239 14949
rect 6181 14940 6193 14943
rect 5500 14912 6193 14940
rect 5500 14900 5506 14912
rect 6181 14909 6193 14912
rect 6227 14909 6239 14943
rect 6181 14903 6239 14909
rect 6638 14900 6644 14952
rect 6696 14900 6702 14952
rect 6730 14900 6736 14952
rect 6788 14940 6794 14952
rect 8220 14940 8248 15116
rect 8570 15036 8576 15088
rect 8628 15076 8634 15088
rect 8757 15079 8815 15085
rect 8757 15076 8769 15079
rect 8628 15048 8769 15076
rect 8628 15036 8634 15048
rect 8757 15045 8769 15048
rect 8803 15045 8815 15079
rect 8757 15039 8815 15045
rect 9493 15079 9551 15085
rect 9493 15045 9505 15079
rect 9539 15076 9551 15079
rect 9766 15076 9772 15088
rect 9539 15048 9772 15076
rect 9539 15045 9551 15048
rect 9493 15039 9551 15045
rect 9766 15036 9772 15048
rect 9824 15036 9830 15088
rect 10134 15036 10140 15088
rect 10192 15036 10198 15088
rect 10796 15076 10824 15116
rect 11882 15104 11888 15156
rect 11940 15104 11946 15156
rect 11977 15147 12035 15153
rect 11977 15113 11989 15147
rect 12023 15144 12035 15147
rect 12158 15144 12164 15156
rect 12023 15116 12164 15144
rect 12023 15113 12035 15116
rect 11977 15107 12035 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12406 15116 13676 15144
rect 12406 15076 12434 15116
rect 10796 15048 12434 15076
rect 12618 15036 12624 15088
rect 12676 15036 12682 15088
rect 13648 15076 13676 15116
rect 13722 15104 13728 15156
rect 13780 15144 13786 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13780 15116 13921 15144
rect 13780 15104 13786 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 16850 15144 16856 15156
rect 13909 15107 13967 15113
rect 14016 15116 16856 15144
rect 14016 15076 14044 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17034 15104 17040 15156
rect 17092 15104 17098 15156
rect 20809 15147 20867 15153
rect 20809 15113 20821 15147
rect 20855 15144 20867 15147
rect 21082 15144 21088 15156
rect 20855 15116 21088 15144
rect 20855 15113 20867 15116
rect 20809 15107 20867 15113
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 13648 15048 14044 15076
rect 15746 15036 15752 15088
rect 15804 15036 15810 15088
rect 16669 15079 16727 15085
rect 16669 15045 16681 15079
rect 16715 15076 16727 15079
rect 17126 15076 17132 15088
rect 16715 15048 17132 15076
rect 16715 15045 16727 15048
rect 16669 15039 16727 15045
rect 17126 15036 17132 15048
rect 17184 15036 17190 15088
rect 10778 14968 10784 15020
rect 10836 15008 10842 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 10836 14980 11713 15008
rect 10836 14968 10842 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 11701 14971 11759 14977
rect 11992 14980 12173 15008
rect 6788 14912 8248 14940
rect 6788 14900 6794 14912
rect 8846 14900 8852 14952
rect 8904 14900 8910 14952
rect 8938 14900 8944 14952
rect 8996 14900 9002 14952
rect 9214 14900 9220 14952
rect 9272 14900 9278 14952
rect 9324 14912 11100 14940
rect 7650 14832 7656 14884
rect 7708 14872 7714 14884
rect 9324 14872 9352 14912
rect 7708 14844 9352 14872
rect 7708 14832 7714 14844
rect 3145 14807 3203 14813
rect 3145 14773 3157 14807
rect 3191 14804 3203 14807
rect 4522 14804 4528 14816
rect 3191 14776 4528 14804
rect 3191 14773 3203 14776
rect 3145 14767 3203 14773
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 8389 14807 8447 14813
rect 8389 14773 8401 14807
rect 8435 14804 8447 14807
rect 9858 14804 9864 14816
rect 8435 14776 9864 14804
rect 8435 14773 8447 14776
rect 8389 14767 8447 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10962 14764 10968 14816
rect 11020 14764 11026 14816
rect 11072 14804 11100 14912
rect 11330 14900 11336 14952
rect 11388 14940 11394 14952
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11388 14912 11529 14940
rect 11388 14900 11394 14912
rect 11517 14909 11529 14912
rect 11563 14940 11575 14943
rect 11790 14940 11796 14952
rect 11563 14912 11796 14940
rect 11563 14909 11575 14912
rect 11517 14903 11575 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 11992 14872 12020 14980
rect 12161 14977 12173 14980
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 12526 14968 12532 15020
rect 12584 14968 12590 15020
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 17310 15008 17316 15020
rect 16899 14980 17316 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 17773 15011 17831 15017
rect 17773 14977 17785 15011
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 12124 14912 14473 14940
rect 12124 14900 12130 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 14734 14900 14740 14952
rect 14792 14900 14798 14952
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 17788 14940 17816 14971
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18693 15011 18751 15017
rect 18693 15008 18705 15011
rect 18104 14980 18705 15008
rect 18104 14968 18110 14980
rect 18693 14977 18705 14980
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 18874 14968 18880 15020
rect 18932 14968 18938 15020
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 20036 14980 20269 15008
rect 20036 14968 20042 14980
rect 20257 14977 20269 14980
rect 20303 15008 20315 15011
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20303 14980 20729 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 18138 14940 18144 14952
rect 16255 14912 18144 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 12618 14872 12624 14884
rect 11992 14844 12624 14872
rect 12618 14832 12624 14844
rect 12676 14832 12682 14884
rect 17865 14875 17923 14881
rect 17865 14841 17877 14875
rect 17911 14872 17923 14875
rect 18322 14872 18328 14884
rect 17911 14844 18328 14872
rect 17911 14841 17923 14844
rect 17865 14835 17923 14841
rect 18322 14832 18328 14844
rect 18380 14832 18386 14884
rect 12250 14804 12256 14816
rect 11072 14776 12256 14804
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 12345 14807 12403 14813
rect 12345 14773 12357 14807
rect 12391 14804 12403 14807
rect 12434 14804 12440 14816
rect 12391 14776 12440 14804
rect 12391 14773 12403 14776
rect 12345 14767 12403 14773
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18141 14807 18199 14813
rect 18141 14804 18153 14807
rect 18012 14776 18153 14804
rect 18012 14764 18018 14776
rect 18141 14773 18153 14776
rect 18187 14773 18199 14807
rect 18141 14767 18199 14773
rect 18506 14764 18512 14816
rect 18564 14804 18570 14816
rect 19061 14807 19119 14813
rect 19061 14804 19073 14807
rect 18564 14776 19073 14804
rect 18564 14764 18570 14776
rect 19061 14773 19073 14776
rect 19107 14773 19119 14807
rect 19061 14767 19119 14773
rect 20070 14764 20076 14816
rect 20128 14764 20134 14816
rect 20254 14764 20260 14816
rect 20312 14804 20318 14816
rect 20349 14807 20407 14813
rect 20349 14804 20361 14807
rect 20312 14776 20361 14804
rect 20312 14764 20318 14776
rect 20349 14773 20361 14776
rect 20395 14773 20407 14807
rect 20349 14767 20407 14773
rect 1104 14714 26312 14736
rect 1104 14662 4101 14714
rect 4153 14662 4165 14714
rect 4217 14662 4229 14714
rect 4281 14662 4293 14714
rect 4345 14662 4357 14714
rect 4409 14662 10403 14714
rect 10455 14662 10467 14714
rect 10519 14662 10531 14714
rect 10583 14662 10595 14714
rect 10647 14662 10659 14714
rect 10711 14662 16705 14714
rect 16757 14662 16769 14714
rect 16821 14662 16833 14714
rect 16885 14662 16897 14714
rect 16949 14662 16961 14714
rect 17013 14662 23007 14714
rect 23059 14662 23071 14714
rect 23123 14662 23135 14714
rect 23187 14662 23199 14714
rect 23251 14662 23263 14714
rect 23315 14662 26312 14714
rect 1104 14640 26312 14662
rect 4890 14560 4896 14612
rect 4948 14560 4954 14612
rect 5718 14560 5724 14612
rect 5776 14560 5782 14612
rect 6365 14603 6423 14609
rect 6365 14569 6377 14603
rect 6411 14600 6423 14603
rect 6638 14600 6644 14612
rect 6411 14572 6644 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 6825 14603 6883 14609
rect 6825 14569 6837 14603
rect 6871 14600 6883 14603
rect 7098 14600 7104 14612
rect 6871 14572 7104 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 11701 14603 11759 14609
rect 11701 14569 11713 14603
rect 11747 14600 11759 14603
rect 12526 14600 12532 14612
rect 11747 14572 12532 14600
rect 11747 14569 11759 14572
rect 11701 14563 11759 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13906 14560 13912 14612
rect 13964 14560 13970 14612
rect 14458 14560 14464 14612
rect 14516 14560 14522 14612
rect 16298 14560 16304 14612
rect 16356 14600 16362 14612
rect 17218 14600 17224 14612
rect 16356 14572 17224 14600
rect 16356 14560 16362 14572
rect 16592 14544 16620 14572
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 18138 14600 18144 14612
rect 17328 14572 18144 14600
rect 6546 14492 6552 14544
rect 6604 14492 6610 14544
rect 8757 14535 8815 14541
rect 8757 14501 8769 14535
rect 8803 14532 8815 14535
rect 11057 14535 11115 14541
rect 8803 14504 9352 14532
rect 8803 14501 8815 14504
rect 8757 14495 8815 14501
rect 6564 14464 6592 14492
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 6564 14436 7021 14464
rect 7009 14433 7021 14436
rect 7055 14464 7067 14467
rect 9214 14464 9220 14476
rect 7055 14436 9220 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9324 14464 9352 14504
rect 11057 14501 11069 14535
rect 11103 14532 11115 14535
rect 11882 14532 11888 14544
rect 11103 14504 11888 14532
rect 11103 14501 11115 14504
rect 11057 14495 11115 14501
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 15194 14532 15200 14544
rect 13464 14504 15200 14532
rect 10870 14464 10876 14476
rect 9324 14436 10876 14464
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11606 14464 11612 14476
rect 11011 14436 11612 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 12124 14436 12173 14464
rect 12124 14424 12130 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12161 14427 12219 14433
rect 12434 14424 12440 14476
rect 12492 14424 12498 14476
rect 12802 14424 12808 14476
rect 12860 14464 12866 14476
rect 13464 14464 13492 14504
rect 15194 14492 15200 14504
rect 15252 14492 15258 14544
rect 16209 14535 16267 14541
rect 16209 14501 16221 14535
rect 16255 14501 16267 14535
rect 16209 14495 16267 14501
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 12860 14436 13492 14464
rect 13556 14436 14657 14464
rect 12860 14424 12866 14436
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4522 14396 4528 14408
rect 4295 14368 4528 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5166 14396 5172 14408
rect 5123 14368 5172 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14396 5687 14399
rect 5994 14396 6000 14408
rect 5675 14368 6000 14396
rect 5675 14365 5687 14368
rect 5629 14359 5687 14365
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 6420 14368 6561 14396
rect 6420 14356 6426 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 6822 14396 6828 14408
rect 6779 14368 6828 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 9122 14356 9128 14408
rect 9180 14356 9186 14408
rect 11241 14399 11299 14405
rect 11241 14365 11253 14399
rect 11287 14365 11299 14399
rect 11241 14359 11299 14365
rect 1946 14288 1952 14340
rect 2004 14328 2010 14340
rect 5534 14328 5540 14340
rect 2004 14300 5540 14328
rect 2004 14288 2010 14300
rect 5534 14288 5540 14300
rect 5592 14328 5598 14340
rect 7285 14331 7343 14337
rect 5592 14300 7236 14328
rect 5592 14288 5598 14300
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 4801 14263 4859 14269
rect 4801 14260 4813 14263
rect 4672 14232 4813 14260
rect 4672 14220 4678 14232
rect 4801 14229 4813 14232
rect 4847 14229 4859 14263
rect 4801 14223 4859 14229
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 6730 14260 6736 14272
rect 5960 14232 6736 14260
rect 5960 14220 5966 14232
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 7208 14260 7236 14300
rect 7285 14297 7297 14331
rect 7331 14328 7343 14331
rect 7374 14328 7380 14340
rect 7331 14300 7380 14328
rect 7331 14297 7343 14300
rect 7285 14291 7343 14297
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 8294 14288 8300 14340
rect 8352 14288 8358 14340
rect 9493 14331 9551 14337
rect 9493 14328 9505 14331
rect 8956 14300 9505 14328
rect 8662 14260 8668 14272
rect 7208 14232 8668 14260
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 8956 14269 8984 14300
rect 9493 14297 9505 14300
rect 9539 14297 9551 14331
rect 9493 14291 9551 14297
rect 10226 14288 10232 14340
rect 10284 14288 10290 14340
rect 8941 14263 8999 14269
rect 8941 14229 8953 14263
rect 8987 14229 8999 14263
rect 11256 14260 11284 14359
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14365 11575 14399
rect 13556 14382 13584 14436
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 16224 14464 16252 14495
rect 16574 14492 16580 14544
rect 16632 14492 16638 14544
rect 17328 14532 17356 14572
rect 18138 14560 18144 14572
rect 18196 14560 18202 14612
rect 17862 14532 17868 14544
rect 16684 14504 17356 14532
rect 17512 14504 17868 14532
rect 16684 14473 16712 14504
rect 14645 14427 14703 14433
rect 15120 14436 16252 14464
rect 16669 14467 16727 14473
rect 11517 14359 11575 14365
rect 11532 14328 11560 14359
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 15120 14405 15148 14436
rect 16669 14433 16681 14467
rect 16715 14433 16727 14467
rect 16669 14427 16727 14433
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14424 14368 14565 14396
rect 14424 14356 14430 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15427 14368 16129 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 16117 14365 16129 14368
rect 16163 14396 16175 14399
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 16163 14368 16497 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 17310 14396 17316 14408
rect 17184 14368 17316 14396
rect 17184 14356 17190 14368
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17512 14405 17540 14504
rect 17862 14492 17868 14504
rect 17920 14532 17926 14544
rect 17920 14504 18874 14532
rect 17920 14492 17926 14504
rect 18233 14467 18291 14473
rect 18233 14433 18245 14467
rect 18279 14464 18291 14467
rect 18279 14436 18736 14464
rect 18279 14433 18291 14436
rect 18233 14427 18291 14433
rect 18708 14408 18736 14436
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 18138 14396 18144 14408
rect 17727 14368 18144 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 12342 14328 12348 14340
rect 11532 14300 12348 14328
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 14093 14331 14151 14337
rect 14093 14297 14105 14331
rect 14139 14297 14151 14331
rect 14093 14291 14151 14297
rect 11514 14260 11520 14272
rect 11256 14232 11520 14260
rect 8941 14223 8999 14229
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14108 14260 14136 14291
rect 14274 14288 14280 14340
rect 14332 14288 14338 14340
rect 14734 14288 14740 14340
rect 14792 14328 14798 14340
rect 14792 14300 15332 14328
rect 14792 14288 14798 14300
rect 13504 14232 14136 14260
rect 13504 14220 13510 14232
rect 15194 14220 15200 14272
rect 15252 14269 15258 14272
rect 15304 14269 15332 14300
rect 15746 14288 15752 14340
rect 15804 14288 15810 14340
rect 15930 14288 15936 14340
rect 15988 14288 15994 14340
rect 16206 14288 16212 14340
rect 16264 14288 16270 14340
rect 17405 14331 17463 14337
rect 17405 14328 17417 14331
rect 16316 14300 17417 14328
rect 15252 14223 15261 14269
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 16316 14260 16344 14300
rect 17405 14297 17417 14300
rect 17451 14297 17463 14331
rect 17405 14291 17463 14297
rect 15335 14232 16344 14260
rect 16393 14263 16451 14269
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 16393 14229 16405 14263
rect 16439 14260 16451 14263
rect 17512 14260 17540 14359
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 18506 14356 18512 14408
rect 18564 14356 18570 14408
rect 18690 14356 18696 14408
rect 18748 14356 18754 14408
rect 18846 14405 18874 14504
rect 19242 14424 19248 14476
rect 19300 14424 19306 14476
rect 18811 14399 18874 14405
rect 18811 14365 18823 14399
rect 18857 14368 18874 14399
rect 18857 14365 18869 14368
rect 18811 14359 18869 14365
rect 18966 14356 18972 14408
rect 19024 14356 19030 14408
rect 18601 14331 18659 14337
rect 18601 14297 18613 14331
rect 18647 14328 18659 14331
rect 19426 14328 19432 14340
rect 18647 14300 19432 14328
rect 18647 14297 18659 14300
rect 18601 14291 18659 14297
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 19521 14331 19579 14337
rect 19521 14297 19533 14331
rect 19567 14297 19579 14331
rect 19521 14291 19579 14297
rect 16439 14232 17540 14260
rect 18325 14263 18383 14269
rect 16439 14229 16451 14232
rect 16393 14223 16451 14229
rect 18325 14229 18337 14263
rect 18371 14260 18383 14263
rect 19536 14260 19564 14291
rect 20070 14288 20076 14340
rect 20128 14288 20134 14340
rect 21269 14331 21327 14337
rect 21269 14297 21281 14331
rect 21315 14297 21327 14331
rect 21269 14291 21327 14297
rect 18371 14232 19564 14260
rect 18371 14229 18383 14232
rect 18325 14223 18383 14229
rect 15252 14220 15258 14223
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 21284 14260 21312 14291
rect 20220 14232 21312 14260
rect 20220 14220 20226 14232
rect 1104 14170 26312 14192
rect 1104 14118 4761 14170
rect 4813 14118 4825 14170
rect 4877 14118 4889 14170
rect 4941 14118 4953 14170
rect 5005 14118 5017 14170
rect 5069 14118 11063 14170
rect 11115 14118 11127 14170
rect 11179 14118 11191 14170
rect 11243 14118 11255 14170
rect 11307 14118 11319 14170
rect 11371 14118 17365 14170
rect 17417 14118 17429 14170
rect 17481 14118 17493 14170
rect 17545 14118 17557 14170
rect 17609 14118 17621 14170
rect 17673 14118 23667 14170
rect 23719 14118 23731 14170
rect 23783 14118 23795 14170
rect 23847 14118 23859 14170
rect 23911 14118 23923 14170
rect 23975 14118 26312 14170
rect 1104 14096 26312 14118
rect 6641 14059 6699 14065
rect 5736 14028 6500 14056
rect 4614 13948 4620 14000
rect 4672 13988 4678 14000
rect 5077 13991 5135 13997
rect 5077 13988 5089 13991
rect 4672 13960 5089 13988
rect 4672 13948 4678 13960
rect 5077 13957 5089 13960
rect 5123 13957 5135 13991
rect 5077 13951 5135 13957
rect 5261 13991 5319 13997
rect 5261 13957 5273 13991
rect 5307 13988 5319 13991
rect 5307 13960 5488 13988
rect 5307 13957 5319 13960
rect 5261 13951 5319 13957
rect 4430 13880 4436 13932
rect 4488 13880 4494 13932
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13889 4767 13923
rect 5460 13920 5488 13960
rect 5736 13929 5764 14028
rect 6472 13988 6500 14028
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 6822 14056 6828 14068
rect 6687 14028 6828 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 7374 14016 7380 14068
rect 7432 14016 7438 14068
rect 8481 14059 8539 14065
rect 8481 14025 8493 14059
rect 8527 14056 8539 14059
rect 9122 14056 9128 14068
rect 8527 14028 9128 14056
rect 8527 14025 8539 14028
rect 8481 14019 8539 14025
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 11149 14059 11207 14065
rect 9548 14028 10916 14056
rect 9548 14016 9554 14028
rect 7466 13988 7472 14000
rect 6472 13960 7472 13988
rect 5721 13923 5779 13929
rect 5460 13892 5672 13920
rect 4709 13883 4767 13889
rect 3878 13812 3884 13864
rect 3936 13852 3942 13864
rect 4724 13852 4752 13883
rect 3936 13824 4752 13852
rect 5644 13852 5672 13892
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 5902 13880 5908 13932
rect 5960 13880 5966 13932
rect 6472 13929 6500 13960
rect 7466 13948 7472 13960
rect 7524 13988 7530 14000
rect 7650 13988 7656 14000
rect 7524 13960 7656 13988
rect 7524 13948 7530 13960
rect 7650 13948 7656 13960
rect 7708 13948 7714 14000
rect 8662 13948 8668 14000
rect 8720 13988 8726 14000
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8720 13960 8861 13988
rect 8720 13948 8726 13960
rect 8849 13957 8861 13960
rect 8895 13957 8907 13991
rect 8849 13951 8907 13957
rect 8941 13991 8999 13997
rect 8941 13957 8953 13991
rect 8987 13988 8999 13991
rect 10042 13988 10048 14000
rect 8987 13960 10048 13988
rect 8987 13957 8999 13960
rect 8941 13951 8999 13957
rect 10042 13948 10048 13960
rect 10100 13948 10106 14000
rect 10778 13948 10784 14000
rect 10836 13948 10842 14000
rect 10888 13988 10916 14028
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11514 14056 11520 14068
rect 11195 14028 11520 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 11790 14056 11796 14068
rect 11624 14028 11796 14056
rect 11624 13988 11652 14028
rect 11790 14016 11796 14028
rect 11848 14056 11854 14068
rect 11974 14056 11980 14068
rect 11848 14028 11980 14056
rect 11848 14016 11854 14028
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 12802 14056 12808 14068
rect 12308 14028 12808 14056
rect 12308 14016 12314 14028
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 12952 14028 13645 14056
rect 12952 14016 12958 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 17126 14016 17132 14068
rect 17184 14056 17190 14068
rect 17494 14056 17500 14068
rect 17184 14028 17500 14056
rect 17184 14016 17190 14028
rect 17494 14016 17500 14028
rect 17552 14056 17558 14068
rect 17957 14059 18015 14065
rect 17957 14056 17969 14059
rect 17552 14028 17969 14056
rect 17552 14016 17558 14028
rect 17957 14025 17969 14028
rect 18003 14025 18015 14059
rect 17957 14019 18015 14025
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18966 14056 18972 14068
rect 18647 14028 18972 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 10888 13960 11652 13988
rect 11882 13948 11888 14000
rect 11940 13988 11946 14000
rect 12161 13991 12219 13997
rect 12161 13988 12173 13991
rect 11940 13960 12173 13988
rect 11940 13948 11946 13960
rect 12161 13957 12173 13960
rect 12207 13957 12219 13991
rect 13817 13991 13875 13997
rect 13817 13988 13829 13991
rect 13386 13960 13829 13988
rect 12161 13951 12219 13957
rect 13817 13957 13829 13960
rect 13863 13957 13875 13991
rect 13817 13951 13875 13957
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 6457 13923 6515 13929
rect 6012 13892 6224 13920
rect 6012 13852 6040 13892
rect 5644 13824 6040 13852
rect 6089 13855 6147 13861
rect 3936 13812 3942 13824
rect 6089 13821 6101 13855
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 4249 13787 4307 13793
rect 4249 13753 4261 13787
rect 4295 13784 4307 13787
rect 6104 13784 6132 13815
rect 4295 13756 6132 13784
rect 6196 13784 6224 13892
rect 6457 13889 6469 13923
rect 6503 13889 6515 13923
rect 6457 13883 6515 13889
rect 7006 13880 7012 13932
rect 7064 13880 7070 13932
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13920 7159 13923
rect 7190 13920 7196 13932
rect 7147 13892 7196 13920
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7190 13880 7196 13892
rect 7248 13880 7254 13932
rect 7282 13880 7288 13932
rect 7340 13920 7346 13932
rect 7561 13923 7619 13929
rect 7561 13920 7573 13923
rect 7340 13892 7573 13920
rect 7340 13880 7346 13892
rect 7561 13889 7573 13892
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 9306 13880 9312 13932
rect 9364 13880 9370 13932
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 10796 13920 10824 13948
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10376 13892 10977 13920
rect 10376 13880 10382 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 13630 13880 13636 13932
rect 13688 13920 13694 13932
rect 13725 13923 13783 13929
rect 13725 13920 13737 13923
rect 13688 13892 13737 13920
rect 13688 13880 13694 13892
rect 13725 13889 13737 13892
rect 13771 13920 13783 13923
rect 14366 13920 14372 13932
rect 13771 13892 14372 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 6730 13784 6736 13796
rect 6196 13756 6736 13784
rect 4295 13753 4307 13756
rect 4249 13747 4307 13753
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 8754 13744 8760 13796
rect 8812 13784 8818 13796
rect 9048 13784 9076 13815
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9548 13824 9597 13852
rect 9548 13812 9554 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 8812 13756 9076 13784
rect 10796 13784 10824 13815
rect 10870 13812 10876 13864
rect 10928 13852 10934 13864
rect 10928 13824 11836 13852
rect 10928 13812 10934 13824
rect 11698 13784 11704 13796
rect 10796 13756 11704 13784
rect 8812 13744 8818 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 11808 13784 11836 13824
rect 11882 13812 11888 13864
rect 11940 13812 11946 13864
rect 14458 13852 14464 13864
rect 11992 13824 14464 13852
rect 11992 13784 12020 13824
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 16298 13852 16304 13864
rect 15804 13824 16304 13852
rect 15804 13812 15810 13824
rect 16298 13812 16304 13824
rect 16356 13852 16362 13864
rect 16942 13852 16948 13864
rect 16356 13824 16948 13852
rect 16356 13812 16362 13824
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 17052 13852 17080 13951
rect 17218 13948 17224 14000
rect 17276 13997 17282 14000
rect 17276 13991 17295 13997
rect 17283 13957 17295 13991
rect 17276 13951 17295 13957
rect 17276 13948 17282 13951
rect 17586 13948 17592 14000
rect 17644 13948 17650 14000
rect 17805 13991 17863 13997
rect 17805 13988 17817 13991
rect 17696 13960 17817 13988
rect 17218 13852 17224 13864
rect 17052 13824 17224 13852
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 11808 13756 12020 13784
rect 17405 13787 17463 13793
rect 17405 13753 17417 13787
rect 17451 13784 17463 13787
rect 17696 13784 17724 13960
rect 17805 13957 17817 13960
rect 17851 13988 17863 13991
rect 18046 13988 18052 14000
rect 17851 13960 18052 13988
rect 17851 13957 17863 13960
rect 17805 13951 17863 13957
rect 18046 13948 18052 13960
rect 18104 13988 18110 14000
rect 18690 13988 18696 14000
rect 18104 13960 18696 13988
rect 18104 13948 18110 13960
rect 18690 13948 18696 13960
rect 18748 13948 18754 14000
rect 20254 13948 20260 14000
rect 20312 13948 20318 14000
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13920 18935 13923
rect 19150 13920 19156 13932
rect 18923 13892 19156 13920
rect 18923 13889 18935 13892
rect 18877 13883 18935 13889
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13821 18199 13855
rect 18141 13815 18199 13821
rect 18248 13852 18276 13883
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 19245 13855 19303 13861
rect 18248 13824 18920 13852
rect 17451 13756 17724 13784
rect 17451 13753 17463 13756
rect 17405 13747 17463 13753
rect 17862 13744 17868 13796
rect 17920 13784 17926 13796
rect 18156 13784 18184 13815
rect 17920 13756 18184 13784
rect 17920 13744 17926 13756
rect 4614 13676 4620 13728
rect 4672 13676 4678 13728
rect 5902 13676 5908 13728
rect 5960 13716 5966 13728
rect 5997 13719 6055 13725
rect 5997 13716 6009 13719
rect 5960 13688 6009 13716
rect 5960 13676 5966 13688
rect 5997 13685 6009 13688
rect 6043 13685 6055 13719
rect 5997 13679 6055 13685
rect 6086 13676 6092 13728
rect 6144 13676 6150 13728
rect 7285 13719 7343 13725
rect 7285 13685 7297 13719
rect 7331 13716 7343 13719
rect 7374 13716 7380 13728
rect 7331 13688 7380 13716
rect 7331 13685 7343 13688
rect 7285 13679 7343 13685
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 11514 13676 11520 13728
rect 11572 13716 11578 13728
rect 11790 13716 11796 13728
rect 11572 13688 11796 13716
rect 11572 13676 11578 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 16482 13676 16488 13728
rect 16540 13716 16546 13728
rect 17221 13719 17279 13725
rect 17221 13716 17233 13719
rect 16540 13688 17233 13716
rect 16540 13676 16546 13688
rect 17221 13685 17233 13688
rect 17267 13685 17279 13719
rect 17221 13679 17279 13685
rect 17773 13719 17831 13725
rect 17773 13685 17785 13719
rect 17819 13716 17831 13719
rect 18248 13716 18276 13824
rect 18892 13796 18920 13824
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19794 13852 19800 13864
rect 19291 13824 19800 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 19794 13812 19800 13824
rect 19852 13812 19858 13864
rect 18874 13744 18880 13796
rect 18932 13744 18938 13796
rect 17819 13688 18276 13716
rect 17819 13685 17831 13688
rect 17773 13679 17831 13685
rect 20346 13676 20352 13728
rect 20404 13716 20410 13728
rect 20671 13719 20729 13725
rect 20671 13716 20683 13719
rect 20404 13688 20683 13716
rect 20404 13676 20410 13688
rect 20671 13685 20683 13688
rect 20717 13685 20729 13719
rect 20671 13679 20729 13685
rect 1104 13626 26312 13648
rect 1104 13574 4101 13626
rect 4153 13574 4165 13626
rect 4217 13574 4229 13626
rect 4281 13574 4293 13626
rect 4345 13574 4357 13626
rect 4409 13574 10403 13626
rect 10455 13574 10467 13626
rect 10519 13574 10531 13626
rect 10583 13574 10595 13626
rect 10647 13574 10659 13626
rect 10711 13574 16705 13626
rect 16757 13574 16769 13626
rect 16821 13574 16833 13626
rect 16885 13574 16897 13626
rect 16949 13574 16961 13626
rect 17013 13574 23007 13626
rect 23059 13574 23071 13626
rect 23123 13574 23135 13626
rect 23187 13574 23199 13626
rect 23251 13574 23263 13626
rect 23315 13574 26312 13626
rect 1104 13552 26312 13574
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 5960 13484 6561 13512
rect 5960 13472 5966 13484
rect 6549 13481 6561 13484
rect 6595 13481 6607 13515
rect 6549 13475 6607 13481
rect 6730 13472 6736 13524
rect 6788 13472 6794 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7101 13515 7159 13521
rect 7101 13512 7113 13515
rect 7064 13484 7113 13512
rect 7064 13472 7070 13484
rect 7101 13481 7113 13484
rect 7147 13512 7159 13515
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 7147 13484 7573 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 7561 13475 7619 13481
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 12618 13512 12624 13524
rect 12575 13484 12624 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 16393 13515 16451 13521
rect 16393 13512 16405 13515
rect 15988 13484 16405 13512
rect 15988 13472 15994 13484
rect 16393 13481 16405 13484
rect 16439 13481 16451 13515
rect 16393 13475 16451 13481
rect 17770 13472 17776 13524
rect 17828 13512 17834 13524
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17828 13484 17877 13512
rect 17828 13472 17834 13484
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18012 13484 19380 13512
rect 18012 13472 18018 13484
rect 5169 13447 5227 13453
rect 5169 13413 5181 13447
rect 5215 13444 5227 13447
rect 5258 13444 5264 13456
rect 5215 13416 5264 13444
rect 5215 13413 5227 13416
rect 5169 13407 5227 13413
rect 5258 13404 5264 13416
rect 5316 13444 5322 13456
rect 5997 13447 6055 13453
rect 5997 13444 6009 13447
rect 5316 13416 6009 13444
rect 5316 13404 5322 13416
rect 5997 13413 6009 13416
rect 6043 13413 6055 13447
rect 5997 13407 6055 13413
rect 7745 13447 7803 13453
rect 7745 13413 7757 13447
rect 7791 13413 7803 13447
rect 7745 13407 7803 13413
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 6086 13376 6092 13388
rect 5399 13348 6092 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 7190 13376 7196 13388
rect 6380 13348 7196 13376
rect 3786 13268 3792 13320
rect 3844 13268 3850 13320
rect 5166 13268 5172 13320
rect 5224 13308 5230 13320
rect 5224 13280 6040 13308
rect 5224 13268 5230 13280
rect 4056 13243 4114 13249
rect 4056 13209 4068 13243
rect 4102 13240 4114 13243
rect 5905 13243 5963 13249
rect 5905 13240 5917 13243
rect 4102 13212 5917 13240
rect 4102 13209 4114 13212
rect 4056 13203 4114 13209
rect 5905 13209 5917 13212
rect 5951 13209 5963 13243
rect 6012 13240 6040 13280
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6380 13317 6408 13348
rect 7190 13336 7196 13348
rect 7248 13376 7254 13388
rect 7760 13376 7788 13407
rect 16298 13404 16304 13456
rect 16356 13404 16362 13456
rect 7248 13348 7788 13376
rect 11333 13379 11391 13385
rect 7248 13336 7254 13348
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11606 13376 11612 13388
rect 11379 13348 11612 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 13446 13376 13452 13388
rect 11716 13348 13452 13376
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6236 13280 6285 13308
rect 6236 13268 6242 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 6656 13240 6684 13271
rect 7650 13268 7656 13320
rect 7708 13268 7714 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10870 13308 10876 13320
rect 10643 13280 10876 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10870 13268 10876 13280
rect 10928 13308 10934 13320
rect 11716 13308 11744 13348
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 15887 13348 16160 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 10928 13280 11744 13308
rect 10928 13268 10934 13280
rect 11790 13268 11796 13320
rect 11848 13308 11854 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 11848 13280 12173 13308
rect 11848 13268 11854 13280
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 12342 13268 12348 13320
rect 12400 13268 12406 13320
rect 12802 13268 12808 13320
rect 12860 13308 12866 13320
rect 13630 13308 13636 13320
rect 12860 13280 13636 13308
rect 12860 13268 12866 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 14090 13268 14096 13320
rect 14148 13268 14154 13320
rect 16022 13268 16028 13320
rect 16080 13268 16086 13320
rect 16132 13317 16160 13348
rect 16868 13348 17325 13376
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 16390 13308 16396 13320
rect 16163 13280 16396 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 6012 13212 6684 13240
rect 7377 13243 7435 13249
rect 5905 13203 5963 13209
rect 7377 13209 7389 13243
rect 7423 13240 7435 13243
rect 7668 13240 7696 13268
rect 7423 13212 7696 13240
rect 7423 13209 7435 13212
rect 7377 13203 7435 13209
rect 10778 13200 10784 13252
rect 10836 13200 10842 13252
rect 10965 13243 11023 13249
rect 10965 13209 10977 13243
rect 11011 13240 11023 13243
rect 12066 13240 12072 13252
rect 11011 13212 12072 13240
rect 11011 13209 11023 13212
rect 10965 13203 11023 13209
rect 12066 13200 12072 13212
rect 12124 13200 12130 13252
rect 14369 13243 14427 13249
rect 14369 13209 14381 13243
rect 14415 13209 14427 13243
rect 14369 13203 14427 13209
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 6181 13175 6239 13181
rect 6181 13172 6193 13175
rect 3568 13144 6193 13172
rect 3568 13132 3574 13144
rect 6181 13141 6193 13144
rect 6227 13141 6239 13175
rect 6181 13135 6239 13141
rect 7282 13132 7288 13184
rect 7340 13172 7346 13184
rect 7577 13175 7635 13181
rect 7577 13172 7589 13175
rect 7340 13144 7589 13172
rect 7340 13132 7346 13144
rect 7577 13141 7589 13144
rect 7623 13141 7635 13175
rect 7577 13135 7635 13141
rect 11514 13132 11520 13184
rect 11572 13172 11578 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11572 13144 11897 13172
rect 11572 13132 11578 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11885 13135 11943 13141
rect 12894 13132 12900 13184
rect 12952 13132 12958 13184
rect 14384 13172 14412 13203
rect 15378 13200 15384 13252
rect 15436 13200 15442 13252
rect 16040 13240 16068 13268
rect 16592 13240 16620 13271
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 16868 13317 16896 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 17788 13376 17816 13472
rect 18141 13447 18199 13453
rect 18141 13413 18153 13447
rect 18187 13444 18199 13447
rect 18874 13444 18880 13456
rect 18187 13416 18880 13444
rect 18187 13413 18199 13416
rect 18141 13407 18199 13413
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 17313 13339 17371 13345
rect 17604 13348 17816 13376
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 17034 13268 17040 13320
rect 17092 13268 17098 13320
rect 17494 13268 17500 13320
rect 17552 13268 17558 13320
rect 16040 13212 16620 13240
rect 16945 13243 17003 13249
rect 16945 13209 16957 13243
rect 16991 13240 17003 13243
rect 17604 13240 17632 13348
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 17920 13348 18245 13376
rect 17920 13336 17926 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18509 13379 18567 13385
rect 18509 13345 18521 13379
rect 18555 13376 18567 13379
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 18555 13348 19257 13376
rect 18555 13345 18567 13348
rect 18509 13339 18567 13345
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 19352 13376 19380 13484
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19852 13484 19901 13512
rect 19852 13472 19858 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 19889 13475 19947 13481
rect 20346 13472 20352 13524
rect 20404 13472 20410 13524
rect 25038 13472 25044 13524
rect 25096 13512 25102 13524
rect 25961 13515 26019 13521
rect 25961 13512 25973 13515
rect 25096 13484 25973 13512
rect 25096 13472 25102 13484
rect 25961 13481 25973 13484
rect 26007 13481 26019 13515
rect 25961 13475 26019 13481
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 20533 13447 20591 13453
rect 20533 13444 20545 13447
rect 19484 13416 20545 13444
rect 19484 13404 19490 13416
rect 20533 13413 20545 13416
rect 20579 13413 20591 13447
rect 20533 13407 20591 13413
rect 19352 13348 20300 13376
rect 19245 13339 19303 13345
rect 17770 13268 17776 13320
rect 17828 13268 17834 13320
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 16991 13212 17632 13240
rect 17681 13243 17739 13249
rect 16991 13209 17003 13212
rect 16945 13203 17003 13209
rect 17681 13209 17693 13243
rect 17727 13240 17739 13243
rect 17954 13240 17960 13252
rect 17727 13212 17960 13240
rect 17727 13209 17739 13212
rect 17681 13203 17739 13209
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 18064 13184 18092 13271
rect 18322 13268 18328 13320
rect 18380 13268 18386 13320
rect 18690 13268 18696 13320
rect 18748 13268 18754 13320
rect 18782 13268 18788 13320
rect 18840 13268 18846 13320
rect 18874 13268 18880 13320
rect 18932 13268 18938 13320
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 15194 13172 15200 13184
rect 14384 13144 15200 13172
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17221 13175 17279 13181
rect 17221 13172 17233 13175
rect 17184 13144 17233 13172
rect 17184 13132 17190 13144
rect 17221 13141 17233 13144
rect 17267 13141 17279 13175
rect 17221 13135 17279 13141
rect 17586 13132 17592 13184
rect 17644 13172 17650 13184
rect 18046 13172 18052 13184
rect 17644 13144 18052 13172
rect 17644 13132 17650 13144
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18598 13132 18604 13184
rect 18656 13172 18662 13184
rect 18984 13172 19012 13271
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19116 13280 19993 13308
rect 19116 13268 19122 13280
rect 19981 13277 19993 13280
rect 20027 13308 20039 13311
rect 20162 13308 20168 13320
rect 20027 13280 20168 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 20272 13317 20300 13348
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 20809 13379 20867 13385
rect 20809 13376 20821 13379
rect 20772 13348 20821 13376
rect 20772 13336 20778 13348
rect 20809 13345 20821 13348
rect 20855 13345 20867 13379
rect 20809 13339 20867 13345
rect 20257 13311 20315 13317
rect 20257 13277 20269 13311
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 25774 13268 25780 13320
rect 25832 13268 25838 13320
rect 21082 13200 21088 13252
rect 21140 13200 21146 13252
rect 23106 13240 23112 13252
rect 22310 13212 23112 13240
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 18656 13144 19012 13172
rect 18656 13132 18662 13144
rect 22370 13132 22376 13184
rect 22428 13172 22434 13184
rect 22557 13175 22615 13181
rect 22557 13172 22569 13175
rect 22428 13144 22569 13172
rect 22428 13132 22434 13144
rect 22557 13141 22569 13144
rect 22603 13141 22615 13175
rect 22557 13135 22615 13141
rect 1104 13082 26312 13104
rect 1104 13030 4761 13082
rect 4813 13030 4825 13082
rect 4877 13030 4889 13082
rect 4941 13030 4953 13082
rect 5005 13030 5017 13082
rect 5069 13030 11063 13082
rect 11115 13030 11127 13082
rect 11179 13030 11191 13082
rect 11243 13030 11255 13082
rect 11307 13030 11319 13082
rect 11371 13030 17365 13082
rect 17417 13030 17429 13082
rect 17481 13030 17493 13082
rect 17545 13030 17557 13082
rect 17609 13030 17621 13082
rect 17673 13030 23667 13082
rect 23719 13030 23731 13082
rect 23783 13030 23795 13082
rect 23847 13030 23859 13082
rect 23911 13030 23923 13082
rect 23975 13030 26312 13082
rect 1104 13008 26312 13030
rect 1504 12940 3464 12968
rect 1504 12909 1532 12940
rect 1489 12903 1547 12909
rect 1489 12869 1501 12903
rect 1535 12869 1547 12903
rect 3436 12900 3464 12940
rect 3510 12928 3516 12980
rect 3568 12928 3574 12980
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 4798 12968 4804 12980
rect 4488 12940 4804 12968
rect 4488 12928 4494 12940
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5166 12928 5172 12980
rect 5224 12928 5230 12980
rect 12802 12968 12808 12980
rect 7024 12940 8248 12968
rect 7024 12900 7052 12940
rect 8220 12900 8248 12940
rect 9692 12940 12808 12968
rect 1489 12863 1547 12869
rect 2148 12872 2774 12900
rect 3436 12872 7052 12900
rect 7116 12872 8064 12900
rect 8220 12872 8708 12900
rect 2148 12776 2176 12872
rect 2222 12792 2228 12844
rect 2280 12832 2286 12844
rect 2389 12835 2447 12841
rect 2389 12832 2401 12835
rect 2280 12804 2401 12832
rect 2280 12792 2286 12804
rect 2389 12801 2401 12804
rect 2435 12801 2447 12835
rect 2746 12832 2774 12872
rect 3786 12832 3792 12844
rect 2746 12804 3792 12832
rect 2389 12795 2447 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4056 12835 4114 12841
rect 4056 12801 4068 12835
rect 4102 12832 4114 12835
rect 4430 12832 4436 12844
rect 4102 12804 4436 12832
rect 4102 12801 4114 12804
rect 4056 12795 4114 12801
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 5258 12792 5264 12844
rect 5316 12792 5322 12844
rect 7116 12841 7144 12872
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12801 7159 12835
rect 7101 12795 7159 12801
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 2130 12724 2136 12776
rect 2188 12724 2194 12776
rect 6457 12767 6515 12773
rect 6457 12733 6469 12767
rect 6503 12764 6515 12767
rect 6546 12764 6552 12776
rect 6503 12736 6552 12764
rect 6503 12733 6515 12736
rect 6457 12727 6515 12733
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 5258 12656 5264 12708
rect 5316 12696 5322 12708
rect 6730 12696 6736 12708
rect 5316 12668 6736 12696
rect 5316 12656 5322 12668
rect 6730 12656 6736 12668
rect 6788 12656 6794 12708
rect 7300 12696 7328 12795
rect 7374 12792 7380 12844
rect 7432 12792 7438 12844
rect 8036 12841 8064 12872
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12832 8079 12835
rect 8570 12832 8576 12844
rect 8067 12804 8576 12832
rect 8067 12801 8079 12804
rect 8021 12795 8079 12801
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 8110 12724 8116 12776
rect 8168 12724 8174 12776
rect 8386 12696 8392 12708
rect 7300 12668 8392 12696
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 8680 12696 8708 12872
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 9692 12832 9720 12940
rect 12802 12928 12808 12940
rect 12860 12968 12866 12980
rect 13078 12968 13084 12980
rect 12860 12940 13084 12968
rect 12860 12928 12866 12940
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 13587 12971 13645 12977
rect 13587 12937 13599 12971
rect 13633 12968 13645 12971
rect 14274 12968 14280 12980
rect 13633 12940 14280 12968
rect 13633 12937 13645 12940
rect 13587 12931 13645 12937
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15378 12928 15384 12980
rect 15436 12928 15442 12980
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12968 16727 12971
rect 17770 12968 17776 12980
rect 16715 12940 17776 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18230 12968 18236 12980
rect 18012 12940 18236 12968
rect 18012 12928 18018 12940
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 18598 12928 18604 12980
rect 18656 12928 18662 12980
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 23106 12928 23112 12980
rect 23164 12928 23170 12980
rect 9950 12860 9956 12912
rect 10008 12900 10014 12912
rect 10008 12872 10456 12900
rect 10008 12860 10014 12872
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9692 12804 9781 12832
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 9858 12792 9864 12844
rect 9916 12792 9922 12844
rect 10042 12792 10048 12844
rect 10100 12792 10106 12844
rect 10134 12792 10140 12844
rect 10192 12792 10198 12844
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 10428 12773 10456 12872
rect 10870 12860 10876 12912
rect 10928 12860 10934 12912
rect 12894 12860 12900 12912
rect 12952 12860 12958 12912
rect 17052 12872 17632 12900
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 8996 12736 10333 12764
rect 8996 12724 9002 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12733 10471 12767
rect 10612 12764 10640 12795
rect 11054 12792 11060 12844
rect 11112 12792 11118 12844
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 11793 12835 11851 12841
rect 11793 12801 11805 12835
rect 11839 12832 11851 12835
rect 11882 12832 11888 12844
rect 11839 12804 11888 12832
rect 11839 12801 11851 12804
rect 11793 12795 11851 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15562 12832 15568 12844
rect 15335 12804 15568 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 16022 12792 16028 12844
rect 16080 12832 16086 12844
rect 17052 12841 17080 12872
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16080 12804 17049 12832
rect 16080 12792 16086 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17310 12792 17316 12844
rect 17368 12792 17374 12844
rect 17604 12841 17632 12872
rect 18046 12860 18052 12912
rect 18104 12900 18110 12912
rect 18104 12872 19104 12900
rect 18104 12860 18110 12872
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12832 18843 12835
rect 18874 12832 18880 12844
rect 18831 12804 18880 12832
rect 18831 12801 18843 12804
rect 18785 12795 18843 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19076 12841 19104 12872
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 20346 12832 20352 12844
rect 19107 12804 20352 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 21232 12804 21373 12832
rect 21232 12792 21238 12804
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 21453 12835 21511 12841
rect 21453 12801 21465 12835
rect 21499 12832 21511 12835
rect 22649 12835 22707 12841
rect 22649 12832 22661 12835
rect 21499 12804 22661 12832
rect 21499 12801 21511 12804
rect 21453 12795 21511 12801
rect 22649 12801 22661 12804
rect 22695 12801 22707 12835
rect 22649 12795 22707 12801
rect 22741 12835 22799 12841
rect 22741 12801 22753 12835
rect 22787 12832 22799 12835
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22787 12804 23029 12832
rect 22787 12801 22799 12804
rect 22741 12795 22799 12801
rect 23017 12801 23029 12804
rect 23063 12832 23075 12835
rect 24670 12832 24676 12844
rect 23063 12804 24676 12832
rect 23063 12801 23075 12804
rect 23017 12795 23075 12801
rect 24670 12792 24676 12804
rect 24728 12792 24734 12844
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 10612 12736 11253 12764
rect 10413 12727 10471 12733
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 9585 12699 9643 12705
rect 8680 12668 8892 12696
rect 1578 12588 1584 12640
rect 1636 12588 1642 12640
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5592 12600 5917 12628
rect 5592 12588 5598 12600
rect 5905 12597 5917 12600
rect 5951 12597 5963 12631
rect 5905 12591 5963 12597
rect 7006 12588 7012 12640
rect 7064 12588 7070 12640
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7466 12628 7472 12640
rect 7147 12600 7472 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 8352 12600 8769 12628
rect 8352 12588 8358 12600
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 8864 12628 8892 12668
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 9674 12696 9680 12708
rect 9631 12668 9680 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 10229 12699 10287 12705
rect 10229 12696 10241 12699
rect 9824 12668 10241 12696
rect 9824 12656 9830 12668
rect 10229 12665 10241 12668
rect 10275 12665 10287 12699
rect 10428 12696 10456 12727
rect 11698 12724 11704 12776
rect 11756 12724 11762 12776
rect 12158 12724 12164 12776
rect 12216 12724 12222 12776
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16540 12736 16865 12764
rect 16540 12724 16546 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17218 12764 17224 12776
rect 17175 12736 17224 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 11716 12696 11744 12724
rect 10428 12668 11744 12696
rect 10229 12659 10287 12665
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 16960 12696 16988 12727
rect 17218 12724 17224 12736
rect 17276 12764 17282 12776
rect 17497 12767 17555 12773
rect 17497 12764 17509 12767
rect 17276 12736 17509 12764
rect 17276 12724 17282 12736
rect 17497 12733 17509 12736
rect 17543 12764 17555 12767
rect 18230 12764 18236 12776
rect 17543 12736 18236 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 21266 12724 21272 12776
rect 21324 12724 21330 12776
rect 21542 12724 21548 12776
rect 21600 12724 21606 12776
rect 22002 12724 22008 12776
rect 22060 12724 22066 12776
rect 16448 12668 17356 12696
rect 16448 12656 16454 12668
rect 10781 12631 10839 12637
rect 10781 12628 10793 12631
rect 8864 12600 10793 12628
rect 8757 12591 8815 12597
rect 10781 12597 10793 12600
rect 10827 12628 10839 12631
rect 11606 12628 11612 12640
rect 10827 12600 11612 12628
rect 10827 12597 10839 12600
rect 10781 12591 10839 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 11701 12631 11759 12637
rect 11701 12597 11713 12631
rect 11747 12628 11759 12631
rect 11790 12628 11796 12640
rect 11747 12600 11796 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 17328 12637 17356 12668
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 18877 12699 18935 12705
rect 18877 12696 18889 12699
rect 18196 12668 18889 12696
rect 18196 12656 18202 12668
rect 18877 12665 18889 12668
rect 18923 12665 18935 12699
rect 18877 12659 18935 12665
rect 18969 12699 19027 12705
rect 18969 12665 18981 12699
rect 19015 12665 19027 12699
rect 18969 12659 19027 12665
rect 17313 12631 17371 12637
rect 17313 12597 17325 12631
rect 17359 12597 17371 12631
rect 17313 12591 17371 12597
rect 17770 12588 17776 12640
rect 17828 12628 17834 12640
rect 18984 12628 19012 12659
rect 17828 12600 19012 12628
rect 17828 12588 17834 12600
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 22833 12631 22891 12637
rect 22833 12628 22845 12631
rect 22336 12600 22845 12628
rect 22336 12588 22342 12600
rect 22833 12597 22845 12600
rect 22879 12597 22891 12631
rect 22833 12591 22891 12597
rect 1104 12538 26312 12560
rect 1104 12486 4101 12538
rect 4153 12486 4165 12538
rect 4217 12486 4229 12538
rect 4281 12486 4293 12538
rect 4345 12486 4357 12538
rect 4409 12486 10403 12538
rect 10455 12486 10467 12538
rect 10519 12486 10531 12538
rect 10583 12486 10595 12538
rect 10647 12486 10659 12538
rect 10711 12486 16705 12538
rect 16757 12486 16769 12538
rect 16821 12486 16833 12538
rect 16885 12486 16897 12538
rect 16949 12486 16961 12538
rect 17013 12486 23007 12538
rect 23059 12486 23071 12538
rect 23123 12486 23135 12538
rect 23187 12486 23199 12538
rect 23251 12486 23263 12538
rect 23315 12486 26312 12538
rect 1104 12464 26312 12486
rect 3050 12424 3056 12436
rect 2056 12396 3056 12424
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12288 1823 12291
rect 2056 12288 2084 12396
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3513 12427 3571 12433
rect 3513 12424 3525 12427
rect 3476 12396 3525 12424
rect 3476 12384 3482 12396
rect 3513 12393 3525 12396
rect 3559 12424 3571 12427
rect 6178 12424 6184 12436
rect 3559 12396 6184 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 7282 12424 7288 12436
rect 6595 12396 7288 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 10965 12427 11023 12433
rect 10965 12393 10977 12427
rect 11011 12424 11023 12427
rect 12158 12424 12164 12436
rect 11011 12396 12164 12424
rect 11011 12393 11023 12396
rect 10965 12387 11023 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 13538 12384 13544 12436
rect 13596 12433 13602 12436
rect 13596 12427 13645 12433
rect 13596 12393 13599 12427
rect 13633 12393 13645 12427
rect 13596 12387 13645 12393
rect 13596 12384 13602 12387
rect 16666 12384 16672 12436
rect 16724 12384 16730 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17129 12427 17187 12433
rect 17129 12424 17141 12427
rect 17092 12396 17141 12424
rect 17092 12384 17098 12396
rect 17129 12393 17141 12396
rect 17175 12393 17187 12427
rect 17129 12387 17187 12393
rect 4798 12316 4804 12368
rect 4856 12356 4862 12368
rect 4856 12328 6316 12356
rect 4856 12316 4862 12328
rect 1811 12260 2084 12288
rect 1811 12257 1823 12260
rect 1765 12251 1823 12257
rect 2130 12248 2136 12300
rect 2188 12248 2194 12300
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 3568 12260 3801 12288
rect 3568 12248 3574 12260
rect 3789 12257 3801 12260
rect 3835 12257 3847 12291
rect 5534 12288 5540 12300
rect 3789 12251 3847 12257
rect 4724 12260 5540 12288
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 3878 12220 3884 12232
rect 1719 12192 3884 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4724 12229 4752 12260
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 6288 12232 6316 12328
rect 8478 12316 8484 12368
rect 8536 12316 8542 12368
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 16531 12359 16589 12365
rect 16531 12356 16543 12359
rect 16448 12328 16543 12356
rect 16448 12316 16454 12328
rect 16531 12325 16543 12328
rect 16577 12325 16589 12359
rect 16684 12356 16712 12384
rect 17310 12356 17316 12368
rect 16684 12328 17316 12356
rect 16531 12319 16589 12325
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6604 12260 7021 12288
rect 6604 12248 6610 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7009 12251 7067 12257
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 10413 12291 10471 12297
rect 8260 12260 8800 12288
rect 8260 12248 8266 12260
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12220 5135 12223
rect 5166 12220 5172 12232
rect 5123 12192 5172 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 6086 12229 6092 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5500 12192 5917 12220
rect 5500 12180 5506 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6053 12223 6092 12229
rect 6053 12189 6065 12223
rect 6053 12183 6092 12189
rect 6086 12180 6092 12183
rect 6144 12180 6150 12232
rect 6270 12180 6276 12232
rect 6328 12180 6334 12232
rect 6370 12223 6428 12229
rect 6370 12189 6382 12223
rect 6416 12189 6428 12223
rect 6370 12183 6428 12189
rect 2400 12155 2458 12161
rect 2400 12121 2412 12155
rect 2446 12152 2458 12155
rect 2498 12152 2504 12164
rect 2446 12124 2504 12152
rect 2446 12121 2458 12124
rect 2400 12115 2458 12121
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 2682 12112 2688 12164
rect 2740 12152 2746 12164
rect 4338 12152 4344 12164
rect 2740 12124 4344 12152
rect 2740 12112 2746 12124
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 5810 12112 5816 12164
rect 5868 12152 5874 12164
rect 6181 12155 6239 12161
rect 6181 12152 6193 12155
rect 5868 12124 6193 12152
rect 5868 12112 5874 12124
rect 6181 12121 6193 12124
rect 6227 12121 6239 12155
rect 6181 12115 6239 12121
rect 2038 12044 2044 12096
rect 2096 12044 2102 12096
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 3844 12056 4445 12084
rect 3844 12044 3850 12056
rect 4433 12053 4445 12056
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 5350 12044 5356 12096
rect 5408 12084 5414 12096
rect 5629 12087 5687 12093
rect 5629 12084 5641 12087
rect 5408 12056 5641 12084
rect 5408 12044 5414 12056
rect 5629 12053 5641 12056
rect 5675 12053 5687 12087
rect 5629 12047 5687 12053
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6385 12084 6413 12183
rect 6638 12180 6644 12232
rect 6696 12180 6702 12232
rect 7276 12223 7334 12229
rect 7276 12189 7288 12223
rect 7322 12220 7334 12223
rect 8294 12220 8300 12232
rect 7322 12192 8300 12220
rect 7322 12189 7334 12192
rect 7276 12183 7334 12189
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12220 8539 12223
rect 8570 12220 8576 12232
rect 8527 12192 8576 12220
rect 8527 12189 8539 12192
rect 8481 12183 8539 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8772 12229 8800 12260
rect 10413 12257 10425 12291
rect 10459 12288 10471 12291
rect 11514 12288 11520 12300
rect 10459 12260 11520 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11747 12260 12173 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 12161 12251 12219 12257
rect 15028 12260 16313 12288
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12220 11207 12223
rect 11606 12220 11612 12232
rect 11195 12192 11612 12220
rect 11195 12189 11207 12192
rect 11149 12183 11207 12189
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 11882 12220 11888 12232
rect 11839 12192 11888 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 8665 12155 8723 12161
rect 8665 12152 8677 12155
rect 6840 12124 8677 12152
rect 6840 12096 6868 12124
rect 8665 12121 8677 12124
rect 8711 12121 8723 12155
rect 8665 12115 8723 12121
rect 9214 12112 9220 12164
rect 9272 12152 9278 12164
rect 11808 12152 11836 12183
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 15028 12229 15056 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12288 16819 12291
rect 16807 12260 17080 12288
rect 16807 12257 16819 12260
rect 16761 12251 16819 12257
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12220 15807 12223
rect 16022 12220 16028 12232
rect 15795 12192 16028 12220
rect 15795 12189 15807 12192
rect 15749 12183 15807 12189
rect 16022 12180 16028 12192
rect 16080 12220 16086 12232
rect 17052 12229 17080 12260
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 22462 12288 22468 12300
rect 21416 12260 22468 12288
rect 21416 12248 21422 12260
rect 22462 12248 22468 12260
rect 22520 12248 22526 12300
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 16080 12192 16405 12220
rect 16080 12180 16086 12192
rect 16393 12189 16405 12192
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17770 12220 17776 12232
rect 17267 12192 17776 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 9272 12124 11836 12152
rect 9272 12112 9278 12124
rect 13170 12112 13176 12164
rect 13228 12112 13234 12164
rect 16868 12152 16896 12183
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 20714 12180 20720 12232
rect 20772 12180 20778 12232
rect 24397 12223 24455 12229
rect 24397 12189 24409 12223
rect 24443 12220 24455 12223
rect 24670 12220 24676 12232
rect 24443 12192 24676 12220
rect 24443 12189 24455 12192
rect 24397 12183 24455 12189
rect 24670 12180 24676 12192
rect 24728 12180 24734 12232
rect 18230 12152 18236 12164
rect 16868 12124 18236 12152
rect 18230 12112 18236 12124
rect 18288 12112 18294 12164
rect 20898 12112 20904 12164
rect 20956 12152 20962 12164
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 20956 12124 21005 12152
rect 20956 12112 20962 12124
rect 20993 12121 21005 12124
rect 21039 12121 21051 12155
rect 22278 12152 22284 12164
rect 22218 12124 22284 12152
rect 20993 12115 21051 12121
rect 22278 12112 22284 12124
rect 22336 12112 22342 12164
rect 22741 12155 22799 12161
rect 22741 12121 22753 12155
rect 22787 12121 22799 12155
rect 22741 12115 22799 12121
rect 6052 12056 6413 12084
rect 6052 12044 6058 12056
rect 6822 12044 6828 12096
rect 6880 12044 6886 12096
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 7708 12056 8401 12084
rect 7708 12044 7714 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8389 12047 8447 12053
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 9640 12056 9965 12084
rect 9640 12044 9646 12056
rect 9953 12053 9965 12056
rect 9999 12053 10011 12087
rect 9953 12047 10011 12053
rect 14550 12044 14556 12096
rect 14608 12084 14614 12096
rect 15105 12087 15163 12093
rect 15105 12084 15117 12087
rect 14608 12056 15117 12084
rect 14608 12044 14614 12056
rect 15105 12053 15117 12056
rect 15151 12053 15163 12087
rect 15105 12047 15163 12053
rect 21174 12044 21180 12096
rect 21232 12084 21238 12096
rect 21910 12084 21916 12096
rect 21232 12056 21916 12084
rect 21232 12044 21238 12056
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 22002 12044 22008 12096
rect 22060 12084 22066 12096
rect 22756 12084 22784 12115
rect 22060 12056 22784 12084
rect 22060 12044 22066 12056
rect 24486 12044 24492 12096
rect 24544 12044 24550 12096
rect 1104 11994 26312 12016
rect 1104 11942 4761 11994
rect 4813 11942 4825 11994
rect 4877 11942 4889 11994
rect 4941 11942 4953 11994
rect 5005 11942 5017 11994
rect 5069 11942 11063 11994
rect 11115 11942 11127 11994
rect 11179 11942 11191 11994
rect 11243 11942 11255 11994
rect 11307 11942 11319 11994
rect 11371 11942 17365 11994
rect 17417 11942 17429 11994
rect 17481 11942 17493 11994
rect 17545 11942 17557 11994
rect 17609 11942 17621 11994
rect 17673 11942 23667 11994
rect 23719 11942 23731 11994
rect 23783 11942 23795 11994
rect 23847 11942 23859 11994
rect 23911 11942 23923 11994
rect 23975 11942 26312 11994
rect 1104 11920 26312 11942
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 2406 11880 2412 11892
rect 2363 11852 2412 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 2406 11840 2412 11852
rect 2464 11880 2470 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2464 11852 2697 11880
rect 2464 11840 2470 11852
rect 2685 11849 2697 11852
rect 2731 11880 2743 11883
rect 2731 11852 3924 11880
rect 2731 11849 2743 11852
rect 2685 11843 2743 11849
rect 2038 11772 2044 11824
rect 2096 11812 2102 11824
rect 2133 11815 2191 11821
rect 2133 11812 2145 11815
rect 2096 11784 2145 11812
rect 2096 11772 2102 11784
rect 2133 11781 2145 11784
rect 2179 11781 2191 11815
rect 2133 11775 2191 11781
rect 2501 11815 2559 11821
rect 2501 11781 2513 11815
rect 2547 11812 2559 11815
rect 2961 11815 3019 11821
rect 2961 11812 2973 11815
rect 2547 11784 2973 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 2961 11781 2973 11784
rect 3007 11781 3019 11815
rect 2961 11775 3019 11781
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2590 11744 2596 11756
rect 2455 11716 2596 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 2884 11676 2912 11707
rect 3050 11704 3056 11756
rect 3108 11704 3114 11756
rect 3234 11704 3240 11756
rect 3292 11704 3298 11756
rect 3418 11704 3424 11756
rect 3476 11704 3482 11756
rect 3786 11704 3792 11756
rect 3844 11704 3850 11756
rect 3896 11744 3924 11852
rect 4338 11840 4344 11892
rect 4396 11840 4402 11892
rect 5810 11840 5816 11892
rect 5868 11840 5874 11892
rect 6086 11840 6092 11892
rect 6144 11880 6150 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 6144 11852 6377 11880
rect 6144 11840 6150 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6638 11840 6644 11892
rect 6696 11880 6702 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 6696 11852 7205 11880
rect 6696 11840 6702 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 7193 11843 7251 11849
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8386 11880 8392 11892
rect 8343 11852 8392 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 9125 11883 9183 11889
rect 9125 11849 9137 11883
rect 9171 11880 9183 11883
rect 10134 11880 10140 11892
rect 9171 11852 10140 11880
rect 9171 11849 9183 11852
rect 9125 11843 9183 11849
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 11011 11883 11069 11889
rect 11011 11880 11023 11883
rect 10836 11852 11023 11880
rect 10836 11840 10842 11852
rect 11011 11849 11023 11852
rect 11057 11849 11069 11883
rect 11011 11843 11069 11849
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11572 11852 11897 11880
rect 11572 11840 11578 11852
rect 11885 11849 11897 11852
rect 11931 11849 11943 11883
rect 11885 11843 11943 11849
rect 13170 11840 13176 11892
rect 13228 11840 13234 11892
rect 14826 11880 14832 11892
rect 14292 11852 14832 11880
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 5534 11812 5540 11824
rect 4028 11784 5540 11812
rect 4028 11772 4034 11784
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 6270 11772 6276 11824
rect 6328 11812 6334 11824
rect 7101 11815 7159 11821
rect 6328 11784 6675 11812
rect 6328 11772 6334 11784
rect 4282 11747 4340 11753
rect 4282 11744 4294 11747
rect 3896 11716 4294 11744
rect 4282 11713 4294 11716
rect 4328 11713 4340 11747
rect 4282 11707 4340 11713
rect 4706 11704 4712 11756
rect 4764 11704 4770 11756
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4948 11716 5181 11744
rect 4948 11704 4954 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5317 11747 5375 11753
rect 5317 11713 5329 11747
rect 5363 11744 5375 11747
rect 5445 11747 5503 11753
rect 5363 11713 5396 11744
rect 5317 11707 5396 11713
rect 5445 11713 5457 11747
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 3605 11679 3663 11685
rect 3605 11676 3617 11679
rect 2884 11648 3617 11676
rect 3605 11645 3617 11648
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 2222 11608 2228 11620
rect 2179 11580 2228 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 2222 11568 2228 11580
rect 2280 11568 2286 11620
rect 2498 11568 2504 11620
rect 2556 11568 2562 11620
rect 3878 11568 3884 11620
rect 3936 11568 3942 11620
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4430 11608 4436 11620
rect 4203 11580 4436 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4430 11568 4436 11580
rect 4488 11568 4494 11620
rect 4816 11540 4844 11639
rect 5368 11608 5396 11707
rect 5460 11676 5488 11707
rect 5631 11704 5637 11756
rect 5689 11704 5695 11756
rect 6086 11704 6092 11756
rect 6144 11744 6150 11756
rect 6380 11744 6500 11754
rect 6647 11753 6675 11784
rect 7101 11781 7113 11815
rect 7147 11812 7159 11815
rect 7374 11812 7380 11824
rect 7147 11784 7380 11812
rect 7147 11781 7159 11784
rect 7101 11775 7159 11781
rect 7374 11772 7380 11784
rect 7432 11772 7438 11824
rect 7561 11815 7619 11821
rect 7561 11781 7573 11815
rect 7607 11812 7619 11815
rect 8110 11812 8116 11824
rect 7607 11784 8116 11812
rect 7607 11781 7619 11784
rect 7561 11775 7619 11781
rect 8110 11772 8116 11784
rect 8168 11772 8174 11824
rect 6532 11747 6590 11753
rect 6532 11744 6544 11747
rect 6144 11742 6316 11744
rect 6380 11742 6544 11744
rect 6144 11726 6544 11742
rect 6144 11716 6408 11726
rect 6472 11716 6544 11726
rect 6144 11704 6150 11716
rect 6288 11714 6408 11716
rect 6532 11713 6544 11716
rect 6578 11713 6590 11747
rect 6532 11707 6590 11713
rect 6642 11747 6700 11753
rect 6642 11713 6654 11747
rect 6688 11713 6700 11747
rect 6642 11707 6700 11713
rect 6730 11704 6736 11756
rect 6788 11742 6794 11756
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6840 11742 6929 11744
rect 6788 11716 6929 11742
rect 6788 11714 6868 11716
rect 6788 11704 6794 11714
rect 6917 11713 6929 11716
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 7466 11704 7472 11756
rect 7524 11704 7530 11756
rect 9582 11704 9588 11756
rect 9640 11704 9646 11756
rect 5994 11676 6000 11688
rect 5460 11648 6000 11676
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 7377 11679 7435 11685
rect 7377 11676 7389 11679
rect 7248 11648 7389 11676
rect 7248 11636 7254 11648
rect 7377 11645 7389 11648
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 7650 11636 7656 11688
rect 7708 11636 7714 11688
rect 8570 11636 8576 11688
rect 8628 11636 8634 11688
rect 9214 11636 9220 11688
rect 9272 11636 9278 11688
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10612 11676 10640 11798
rect 11164 11784 12434 11812
rect 11164 11753 11192 11784
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 11974 11744 11980 11756
rect 11931 11716 11980 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 10100 11648 10548 11676
rect 10612 11648 11253 11676
rect 10100 11636 10106 11648
rect 6270 11608 6276 11620
rect 5368 11580 6276 11608
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 10520 11608 10548 11648
rect 11241 11645 11253 11648
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 10962 11608 10968 11620
rect 10520 11580 10968 11608
rect 10962 11568 10968 11580
rect 11020 11608 11026 11620
rect 11532 11608 11560 11707
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 12124 11716 12173 11744
rect 12124 11704 12130 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12406 11744 12434 11784
rect 13078 11744 13084 11756
rect 12406 11716 13084 11744
rect 12161 11707 12219 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14292 11753 14320 11852
rect 14826 11840 14832 11852
rect 14884 11880 14890 11892
rect 14884 11852 16712 11880
rect 14884 11840 14890 11852
rect 14550 11772 14556 11824
rect 14608 11772 14614 11824
rect 16301 11815 16359 11821
rect 16301 11812 16313 11815
rect 15778 11784 16313 11812
rect 16301 11781 16313 11784
rect 16347 11781 16359 11815
rect 16301 11775 16359 11781
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 14148 11716 14289 11744
rect 14148 11704 14154 11716
rect 14277 11713 14289 11716
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16684 11744 16712 11852
rect 18782 11840 18788 11892
rect 18840 11889 18846 11892
rect 18840 11883 18859 11889
rect 18847 11849 18859 11883
rect 18840 11843 18859 11849
rect 18840 11840 18846 11843
rect 20898 11840 20904 11892
rect 20956 11840 20962 11892
rect 21450 11880 21456 11892
rect 21008 11852 21456 11880
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 17126 11812 17132 11824
rect 17083 11784 17132 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 17126 11772 17132 11784
rect 17184 11772 17190 11824
rect 17770 11772 17776 11824
rect 17828 11772 17834 11824
rect 18414 11772 18420 11824
rect 18472 11812 18478 11824
rect 18601 11815 18659 11821
rect 18601 11812 18613 11815
rect 18472 11784 18613 11812
rect 18472 11772 18478 11784
rect 18601 11781 18613 11784
rect 18647 11781 18659 11815
rect 21008 11812 21036 11852
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21600 11852 21833 11880
rect 21600 11840 21606 11852
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 23474 11880 23480 11892
rect 21821 11843 21879 11849
rect 22066 11852 23480 11880
rect 18601 11775 18659 11781
rect 20916 11784 21036 11812
rect 21100 11784 21680 11812
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 16684 11716 16773 11744
rect 16209 11707 16267 11713
rect 16761 11713 16773 11716
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 20441 11747 20499 11753
rect 20441 11713 20453 11747
rect 20487 11744 20499 11747
rect 20806 11744 20812 11756
rect 20487 11716 20812 11744
rect 20487 11713 20499 11716
rect 20441 11707 20499 11713
rect 11790 11636 11796 11688
rect 11848 11636 11854 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12986 11676 12992 11688
rect 12483 11648 12992 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 12986 11636 12992 11648
rect 13044 11636 13050 11688
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 16224 11676 16252 11707
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 18322 11676 18328 11688
rect 15620 11648 16252 11676
rect 16868 11648 18328 11676
rect 15620 11636 15626 11648
rect 12158 11608 12164 11620
rect 11020 11580 12164 11608
rect 11020 11568 11026 11580
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 15654 11568 15660 11620
rect 15712 11608 15718 11620
rect 16868 11608 16896 11648
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11676 20591 11679
rect 20916 11676 20944 11784
rect 21100 11753 21128 11784
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 21174 11704 21180 11756
rect 21232 11704 21238 11756
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11713 21327 11747
rect 21269 11707 21327 11713
rect 20579 11648 20944 11676
rect 20579 11645 20591 11648
rect 20533 11639 20591 11645
rect 20990 11636 20996 11688
rect 21048 11676 21054 11688
rect 21284 11676 21312 11707
rect 21358 11704 21364 11756
rect 21416 11753 21422 11756
rect 21416 11747 21445 11753
rect 21433 11713 21445 11747
rect 21416 11707 21445 11713
rect 21416 11704 21422 11707
rect 21048 11648 21312 11676
rect 21545 11679 21603 11685
rect 21048 11636 21054 11648
rect 21545 11645 21557 11679
rect 21591 11645 21603 11679
rect 21652 11676 21680 11784
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 22066 11812 22094 11852
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 24492 11824 24544 11830
rect 21968 11784 22140 11812
rect 21968 11772 21974 11784
rect 21818 11704 21824 11756
rect 21876 11744 21882 11756
rect 22002 11744 22008 11756
rect 21876 11716 22008 11744
rect 21876 11704 21882 11716
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22112 11753 22140 11784
rect 22186 11772 22192 11824
rect 22244 11812 22250 11824
rect 22649 11815 22707 11821
rect 22649 11812 22661 11815
rect 22244 11784 22661 11812
rect 22244 11772 22250 11784
rect 22649 11781 22661 11784
rect 22695 11781 22707 11815
rect 22649 11775 22707 11781
rect 24492 11766 24544 11772
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22370 11744 22376 11756
rect 22327 11716 22376 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 22462 11704 22468 11756
rect 22520 11744 22526 11756
rect 22922 11744 22928 11756
rect 22520 11716 22928 11744
rect 22520 11704 22526 11716
rect 22922 11704 22928 11716
rect 22980 11704 22986 11756
rect 23106 11704 23112 11756
rect 23164 11704 23170 11756
rect 24578 11704 24584 11756
rect 24636 11744 24642 11756
rect 24949 11747 25007 11753
rect 24949 11744 24961 11747
rect 24636 11716 24961 11744
rect 24636 11704 24642 11716
rect 24949 11713 24961 11716
rect 24995 11744 25007 11747
rect 25041 11747 25099 11753
rect 25041 11744 25053 11747
rect 24995 11716 25053 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 25041 11713 25053 11716
rect 25087 11713 25099 11747
rect 25041 11707 25099 11713
rect 22833 11679 22891 11685
rect 22833 11676 22845 11679
rect 21652 11648 22845 11676
rect 21545 11639 21603 11645
rect 22833 11645 22845 11648
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 23477 11679 23535 11685
rect 23477 11645 23489 11679
rect 23523 11676 23535 11679
rect 24026 11676 24032 11688
rect 23523 11648 24032 11676
rect 23523 11645 23535 11648
rect 23477 11639 23535 11645
rect 15712 11580 16896 11608
rect 18340 11608 18368 11636
rect 20809 11611 20867 11617
rect 18340 11580 18828 11608
rect 15712 11568 15718 11580
rect 5902 11540 5908 11552
rect 4816 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 11609 11543 11667 11549
rect 11609 11540 11621 11543
rect 11572 11512 11621 11540
rect 11572 11500 11578 11512
rect 11609 11509 11621 11512
rect 11655 11509 11667 11543
rect 11609 11503 11667 11509
rect 16022 11500 16028 11552
rect 16080 11500 16086 11552
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18800 11549 18828 11580
rect 20809 11577 20821 11611
rect 20855 11608 20867 11611
rect 21560 11608 21588 11639
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 20855 11580 21588 11608
rect 20855 11577 20867 11580
rect 20809 11571 20867 11577
rect 21634 11568 21640 11620
rect 21692 11608 21698 11620
rect 22189 11611 22247 11617
rect 22189 11608 22201 11611
rect 21692 11580 22201 11608
rect 21692 11568 21698 11580
rect 22189 11577 22201 11580
rect 22235 11577 22247 11611
rect 24946 11608 24952 11620
rect 22189 11571 22247 11577
rect 24780 11580 24952 11608
rect 18509 11543 18567 11549
rect 18509 11540 18521 11543
rect 18288 11512 18521 11540
rect 18288 11500 18294 11512
rect 18509 11509 18521 11512
rect 18555 11509 18567 11543
rect 18509 11503 18567 11509
rect 18785 11543 18843 11549
rect 18785 11509 18797 11543
rect 18831 11509 18843 11543
rect 18785 11503 18843 11509
rect 18969 11543 19027 11549
rect 18969 11509 18981 11543
rect 19015 11540 19027 11543
rect 19426 11540 19432 11552
rect 19015 11512 19432 11540
rect 19015 11509 19027 11512
rect 18969 11503 19027 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 20898 11500 20904 11552
rect 20956 11540 20962 11552
rect 21450 11540 21456 11552
rect 20956 11512 21456 11540
rect 20956 11500 20962 11512
rect 21450 11500 21456 11512
rect 21508 11540 21514 11552
rect 21818 11540 21824 11552
rect 21508 11512 21824 11540
rect 21508 11500 21514 11512
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 22002 11500 22008 11552
rect 22060 11540 22066 11552
rect 23934 11540 23940 11552
rect 22060 11512 23940 11540
rect 22060 11500 22066 11512
rect 23934 11500 23940 11512
rect 23992 11540 23998 11552
rect 24780 11540 24808 11580
rect 24946 11568 24952 11580
rect 25004 11568 25010 11620
rect 23992 11512 24808 11540
rect 23992 11500 23998 11512
rect 25682 11500 25688 11552
rect 25740 11500 25746 11552
rect 1104 11450 26312 11472
rect 1104 11398 4101 11450
rect 4153 11398 4165 11450
rect 4217 11398 4229 11450
rect 4281 11398 4293 11450
rect 4345 11398 4357 11450
rect 4409 11398 10403 11450
rect 10455 11398 10467 11450
rect 10519 11398 10531 11450
rect 10583 11398 10595 11450
rect 10647 11398 10659 11450
rect 10711 11398 16705 11450
rect 16757 11398 16769 11450
rect 16821 11398 16833 11450
rect 16885 11398 16897 11450
rect 16949 11398 16961 11450
rect 17013 11398 23007 11450
rect 23059 11398 23071 11450
rect 23123 11398 23135 11450
rect 23187 11398 23199 11450
rect 23251 11398 23263 11450
rect 23315 11398 26312 11450
rect 1104 11376 26312 11398
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3881 11339 3939 11345
rect 3881 11336 3893 11339
rect 3108 11308 3893 11336
rect 3108 11296 3114 11308
rect 3881 11305 3893 11308
rect 3927 11336 3939 11339
rect 4614 11336 4620 11348
rect 3927 11308 4620 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 4890 11296 4896 11348
rect 4948 11296 4954 11348
rect 5000 11308 5396 11336
rect 3326 11228 3332 11280
rect 3384 11268 3390 11280
rect 4709 11271 4767 11277
rect 4709 11268 4721 11271
rect 3384 11240 4721 11268
rect 3384 11228 3390 11240
rect 4709 11237 4721 11240
rect 4755 11268 4767 11271
rect 5000 11268 5028 11308
rect 4755 11240 5028 11268
rect 4755 11237 4767 11240
rect 4709 11231 4767 11237
rect 5258 11228 5264 11280
rect 5316 11228 5322 11280
rect 5368 11268 5396 11308
rect 5442 11296 5448 11348
rect 5500 11296 5506 11348
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 5552 11308 5641 11336
rect 5552 11280 5580 11308
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 5629 11299 5687 11305
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 6328 11308 6561 11336
rect 6328 11296 6334 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8628 11308 8769 11336
rect 8628 11296 8634 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 11054 11345 11060 11348
rect 11011 11339 11060 11345
rect 8904 11308 10916 11336
rect 8904 11296 8910 11308
rect 5534 11268 5540 11280
rect 5368 11240 5540 11268
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 5718 11228 5724 11280
rect 5776 11268 5782 11280
rect 6362 11268 6368 11280
rect 5776 11240 6368 11268
rect 5776 11228 5782 11240
rect 6362 11228 6368 11240
rect 6420 11228 6426 11280
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11200 5043 11203
rect 5166 11200 5172 11212
rect 5031 11172 5172 11200
rect 5031 11169 5043 11172
rect 4985 11163 5043 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6270 11200 6276 11212
rect 6135 11172 6276 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 7190 11200 7196 11212
rect 6380 11172 7196 11200
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3292 11104 3801 11132
rect 3292 11092 3298 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4019 11104 4445 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4433 11101 4445 11104
rect 4479 11132 4491 11135
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 4479 11104 5549 11132
rect 4479 11101 4491 11104
rect 4433 11095 4491 11101
rect 5537 11101 5549 11104
rect 5583 11132 5595 11135
rect 6178 11132 6184 11144
rect 5583 11104 6184 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 3804 11064 3832 11095
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6380 11064 6408 11172
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 9585 11203 9643 11209
rect 9585 11169 9597 11203
rect 9631 11200 9643 11203
rect 9766 11200 9772 11212
rect 9631 11172 9772 11200
rect 9631 11169 9643 11172
rect 9585 11163 9643 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 6604 11104 7389 11132
rect 6604 11092 6610 11104
rect 7377 11101 7389 11104
rect 7423 11132 7435 11135
rect 9214 11132 9220 11144
rect 7423 11104 9220 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 3804 11036 6408 11064
rect 6454 11024 6460 11076
rect 6512 11064 6518 11076
rect 6733 11067 6791 11073
rect 6733 11064 6745 11067
rect 6512 11036 6745 11064
rect 6512 11024 6518 11036
rect 6733 11033 6745 11036
rect 6779 11033 6791 11067
rect 6733 11027 6791 11033
rect 7644 11067 7702 11073
rect 7644 11033 7656 11067
rect 7690 11064 7702 11067
rect 8478 11064 8484 11076
rect 7690 11036 8484 11064
rect 7690 11033 7702 11036
rect 7644 11027 7702 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9950 11024 9956 11076
rect 10008 11024 10014 11076
rect 10888 11064 10916 11308
rect 11011 11305 11023 11339
rect 11057 11305 11060 11339
rect 11011 11299 11060 11305
rect 11054 11296 11060 11299
rect 11112 11296 11118 11348
rect 11606 11296 11612 11348
rect 11664 11296 11670 11348
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 11848 11308 12112 11336
rect 11848 11296 11854 11308
rect 11333 11271 11391 11277
rect 11333 11237 11345 11271
rect 11379 11268 11391 11271
rect 11974 11268 11980 11280
rect 11379 11240 11980 11268
rect 11379 11237 11391 11240
rect 11333 11231 11391 11237
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 11698 11200 11704 11212
rect 11655 11172 11704 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 12084 11200 12112 11308
rect 12158 11296 12164 11348
rect 12216 11296 12222 11348
rect 15654 11336 15660 11348
rect 13648 11308 15660 11336
rect 11808 11172 12434 11200
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11241 11135 11299 11141
rect 11241 11132 11253 11135
rect 11020 11104 11253 11132
rect 11020 11092 11026 11104
rect 11241 11101 11253 11104
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11132 11575 11135
rect 11808 11132 11836 11172
rect 12406 11144 12434 11172
rect 11563 11104 11836 11132
rect 11563 11101 11575 11104
rect 11517 11095 11575 11101
rect 11882 11092 11888 11144
rect 11940 11092 11946 11144
rect 12406 11104 12440 11144
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 11698 11064 11704 11076
rect 10888 11036 11704 11064
rect 11698 11024 11704 11036
rect 11756 11064 11762 11076
rect 13648 11064 13676 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 15764 11308 16712 11336
rect 15764 11268 15792 11308
rect 14200 11240 15792 11268
rect 15841 11271 15899 11277
rect 14200 11200 14228 11240
rect 15841 11237 15853 11271
rect 15887 11268 15899 11271
rect 16574 11268 16580 11280
rect 15887 11240 16580 11268
rect 15887 11237 15899 11240
rect 15841 11231 15899 11237
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 16684 11268 16712 11308
rect 17770 11296 17776 11348
rect 17828 11336 17834 11348
rect 17865 11339 17923 11345
rect 17865 11336 17877 11339
rect 17828 11308 17877 11336
rect 17828 11296 17834 11308
rect 17865 11305 17877 11308
rect 17911 11305 17923 11339
rect 20806 11336 20812 11348
rect 17865 11299 17923 11305
rect 19812 11308 20812 11336
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 16684 11240 19257 11268
rect 19245 11237 19257 11240
rect 19291 11237 19303 11271
rect 19245 11231 19303 11237
rect 17954 11200 17960 11212
rect 13740 11172 14228 11200
rect 13740 11141 13768 11172
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14200 11141 14228 11172
rect 14844 11172 17960 11200
rect 14844 11141 14872 11172
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18046 11160 18052 11212
rect 18104 11200 18110 11212
rect 18233 11203 18291 11209
rect 18233 11200 18245 11203
rect 18104 11172 18245 11200
rect 18104 11160 18110 11172
rect 18233 11169 18245 11172
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 18322 11160 18328 11212
rect 18380 11160 18386 11212
rect 19702 11160 19708 11212
rect 19760 11160 19766 11212
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 13872 11104 13921 11132
rect 13872 11092 13878 11104
rect 13909 11101 13921 11104
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 14185 11135 14243 11141
rect 14185 11101 14197 11135
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 14829 11135 14887 11141
rect 14829 11132 14841 11135
rect 14599 11104 14841 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 14829 11101 14841 11104
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 11756 11036 13676 11064
rect 13924 11064 13952 11095
rect 15010 11092 15016 11144
rect 15068 11092 15074 11144
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 15620 11104 17785 11132
rect 15620 11092 15626 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 19812 11141 19840 11308
rect 20806 11296 20812 11308
rect 20864 11336 20870 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20864 11308 20913 11336
rect 20864 11296 20870 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 21913 11339 21971 11345
rect 21913 11336 21925 11339
rect 20901 11299 20959 11305
rect 21008 11308 21925 11336
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11101 19855 11135
rect 21008 11132 21036 11308
rect 21913 11305 21925 11308
rect 21959 11336 21971 11339
rect 22278 11336 22284 11348
rect 21959 11308 22284 11336
rect 21959 11305 21971 11308
rect 21913 11299 21971 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22833 11339 22891 11345
rect 22833 11336 22845 11339
rect 22572 11308 22845 11336
rect 21085 11271 21143 11277
rect 21085 11237 21097 11271
rect 21131 11237 21143 11271
rect 21085 11231 21143 11237
rect 21100 11200 21128 11231
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 22373 11271 22431 11277
rect 22373 11268 22385 11271
rect 21232 11240 22385 11268
rect 21232 11228 21238 11240
rect 22373 11237 22385 11240
rect 22419 11237 22431 11271
rect 22373 11231 22431 11237
rect 22002 11200 22008 11212
rect 21100 11172 22008 11200
rect 22002 11160 22008 11172
rect 22060 11160 22066 11212
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11200 22155 11203
rect 22186 11200 22192 11212
rect 22143 11172 22192 11200
rect 22143 11169 22155 11172
rect 22097 11163 22155 11169
rect 22186 11160 22192 11172
rect 22244 11200 22250 11212
rect 22572 11200 22600 11308
rect 22833 11305 22845 11308
rect 22879 11305 22891 11339
rect 24026 11336 24032 11348
rect 22833 11299 22891 11305
rect 23768 11308 24032 11336
rect 23566 11228 23572 11280
rect 23624 11268 23630 11280
rect 23661 11271 23719 11277
rect 23661 11268 23673 11271
rect 23624 11240 23673 11268
rect 23624 11228 23630 11240
rect 23661 11237 23673 11240
rect 23707 11237 23719 11271
rect 23661 11231 23719 11237
rect 23474 11200 23480 11212
rect 22244 11172 22600 11200
rect 22664 11172 23480 11200
rect 22244 11160 22250 11172
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 19797 11095 19855 11101
rect 20732 11104 21373 11132
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 13924 11036 14381 11064
rect 11756 11024 11762 11036
rect 14369 11033 14381 11036
rect 14415 11033 14427 11067
rect 14369 11027 14427 11033
rect 14461 11067 14519 11073
rect 14461 11033 14473 11067
rect 14507 11064 14519 11067
rect 15028 11064 15056 11092
rect 14507 11036 15056 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 15470 11024 15476 11076
rect 15528 11064 15534 11076
rect 15689 11067 15747 11073
rect 15528 11036 15608 11064
rect 15528 11024 15534 11036
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 5258 10996 5264 11008
rect 4488 10968 5264 10996
rect 4488 10956 4494 10968
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 6086 10956 6092 11008
rect 6144 10996 6150 11008
rect 6825 10999 6883 11005
rect 6825 10996 6837 10999
rect 6144 10968 6837 10996
rect 6144 10956 6150 10968
rect 6825 10965 6837 10968
rect 6871 10965 6883 10999
rect 6825 10959 6883 10965
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 13817 10999 13875 11005
rect 13817 10996 13829 10999
rect 13688 10968 13829 10996
rect 13688 10956 13694 10968
rect 13817 10965 13829 10968
rect 13863 10965 13875 10999
rect 13817 10959 13875 10965
rect 14734 10956 14740 11008
rect 14792 10956 14798 11008
rect 14918 10956 14924 11008
rect 14976 10956 14982 11008
rect 15580 10996 15608 11036
rect 15689 11033 15701 11067
rect 15735 11064 15747 11067
rect 16022 11064 16028 11076
rect 15735 11036 16028 11064
rect 15735 11033 15747 11036
rect 15689 11027 15747 11033
rect 16022 11024 16028 11036
rect 16080 11024 16086 11076
rect 17034 11064 17040 11076
rect 16132 11036 17040 11064
rect 16132 10996 16160 11036
rect 17034 11024 17040 11036
rect 17092 11064 17098 11076
rect 18432 11064 18460 11092
rect 17092 11036 18460 11064
rect 17092 11024 17098 11036
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 19536 11064 19564 11095
rect 20732 11073 20760 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 21450 11092 21456 11144
rect 21508 11092 21514 11144
rect 21542 11092 21548 11144
rect 21600 11092 21606 11144
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11134 21695 11135
rect 21683 11106 21772 11134
rect 21683 11101 21695 11106
rect 21637 11095 21695 11101
rect 20717 11067 20775 11073
rect 20717 11064 20729 11067
rect 18748 11036 19564 11064
rect 20640 11036 20729 11064
rect 18748 11024 18754 11036
rect 15580 10968 16160 10996
rect 18049 10999 18107 11005
rect 18049 10965 18061 10999
rect 18095 10996 18107 10999
rect 18414 10996 18420 11008
rect 18095 10968 18420 10996
rect 18095 10965 18107 10968
rect 18049 10959 18107 10965
rect 18414 10956 18420 10968
rect 18472 10956 18478 11008
rect 18782 10956 18788 11008
rect 18840 10996 18846 11008
rect 20640 10996 20668 11036
rect 20717 11033 20729 11036
rect 20763 11033 20775 11067
rect 20717 11027 20775 11033
rect 20933 11067 20991 11073
rect 20933 11033 20945 11067
rect 20979 11064 20991 11067
rect 21266 11064 21272 11076
rect 20979 11036 21272 11064
rect 20979 11033 20991 11036
rect 20933 11027 20991 11033
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 21744 11064 21772 11106
rect 21818 11092 21824 11144
rect 21876 11092 21882 11144
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11132 22523 11135
rect 22664 11132 22692 11172
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 23768 11200 23796 11308
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24397 11271 24455 11277
rect 24397 11268 24409 11271
rect 23584 11172 23796 11200
rect 23860 11240 24409 11268
rect 22511 11104 22692 11132
rect 22741 11135 22799 11141
rect 22511 11101 22523 11104
rect 22465 11095 22523 11101
rect 22741 11101 22753 11135
rect 22787 11132 22799 11135
rect 22922 11132 22928 11144
rect 22787 11104 22928 11132
rect 22787 11101 22799 11104
rect 22741 11095 22799 11101
rect 22922 11092 22928 11104
rect 22980 11092 22986 11144
rect 22557 11067 22615 11073
rect 22557 11064 22569 11067
rect 21744 11036 22569 11064
rect 22557 11033 22569 11036
rect 22603 11033 22615 11067
rect 23584 11064 23612 11172
rect 23661 11135 23719 11141
rect 23661 11101 23673 11135
rect 23707 11132 23719 11135
rect 23860 11132 23888 11240
rect 24397 11237 24409 11240
rect 24443 11237 24455 11271
rect 24397 11231 24455 11237
rect 25682 11200 25688 11212
rect 24412 11172 25688 11200
rect 23707 11104 23888 11132
rect 23937 11135 23995 11141
rect 23707 11101 23719 11104
rect 23661 11095 23719 11101
rect 23937 11101 23949 11135
rect 23983 11101 23995 11135
rect 23937 11095 23995 11101
rect 23845 11067 23903 11073
rect 23845 11064 23857 11067
rect 22557 11027 22615 11033
rect 22664 11036 23520 11064
rect 23584 11036 23857 11064
rect 18840 10968 20668 10996
rect 21177 10999 21235 11005
rect 18840 10956 18846 10968
rect 21177 10965 21189 10999
rect 21223 10996 21235 10999
rect 21358 10996 21364 11008
rect 21223 10968 21364 10996
rect 21223 10965 21235 10968
rect 21177 10959 21235 10965
rect 21358 10956 21364 10968
rect 21416 10996 21422 11008
rect 22664 10996 22692 11036
rect 21416 10968 22692 10996
rect 23492 10996 23520 11036
rect 23845 11033 23857 11036
rect 23891 11033 23903 11067
rect 23952 11064 23980 11095
rect 24026 11092 24032 11144
rect 24084 11092 24090 11144
rect 24210 11092 24216 11144
rect 24268 11092 24274 11144
rect 24412 11141 24440 11172
rect 25682 11160 25688 11172
rect 25740 11160 25746 11212
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24673 11135 24731 11141
rect 24673 11101 24685 11135
rect 24719 11101 24731 11135
rect 24673 11095 24731 11101
rect 24118 11064 24124 11076
rect 23952 11036 24124 11064
rect 23845 11027 23903 11033
rect 24118 11024 24124 11036
rect 24176 11064 24182 11076
rect 24688 11064 24716 11095
rect 24176 11036 24716 11064
rect 24176 11024 24182 11036
rect 24210 10996 24216 11008
rect 23492 10968 24216 10996
rect 21416 10956 21422 10968
rect 24210 10956 24216 10968
rect 24268 10996 24274 11008
rect 24581 10999 24639 11005
rect 24581 10996 24593 10999
rect 24268 10968 24593 10996
rect 24268 10956 24274 10968
rect 24581 10965 24593 10968
rect 24627 10965 24639 10999
rect 24581 10959 24639 10965
rect 1104 10906 26312 10928
rect 1104 10854 4761 10906
rect 4813 10854 4825 10906
rect 4877 10854 4889 10906
rect 4941 10854 4953 10906
rect 5005 10854 5017 10906
rect 5069 10854 11063 10906
rect 11115 10854 11127 10906
rect 11179 10854 11191 10906
rect 11243 10854 11255 10906
rect 11307 10854 11319 10906
rect 11371 10854 17365 10906
rect 17417 10854 17429 10906
rect 17481 10854 17493 10906
rect 17545 10854 17557 10906
rect 17609 10854 17621 10906
rect 17673 10854 23667 10906
rect 23719 10854 23731 10906
rect 23783 10854 23795 10906
rect 23847 10854 23859 10906
rect 23911 10854 23923 10906
rect 23975 10854 26312 10906
rect 1104 10832 26312 10854
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6565 10795 6623 10801
rect 6565 10792 6577 10795
rect 5500 10764 6577 10792
rect 5500 10752 5506 10764
rect 6565 10761 6577 10764
rect 6611 10761 6623 10795
rect 6565 10755 6623 10761
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9306 10792 9312 10804
rect 9171 10764 9312 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 11698 10752 11704 10804
rect 11756 10752 11762 10804
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18012 10764 18245 10792
rect 18012 10752 18018 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 18322 10752 18328 10804
rect 18380 10792 18386 10804
rect 18380 10764 19380 10792
rect 18380 10752 18386 10764
rect 2406 10684 2412 10736
rect 2464 10684 2470 10736
rect 2625 10727 2683 10733
rect 2625 10693 2637 10727
rect 2671 10724 2683 10727
rect 2866 10724 2872 10736
rect 2671 10696 2872 10724
rect 2671 10693 2683 10696
rect 2625 10687 2683 10693
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 19352 10733 19380 10764
rect 22186 10752 22192 10804
rect 22244 10752 22250 10804
rect 24029 10795 24087 10801
rect 24029 10761 24041 10795
rect 24075 10792 24087 10795
rect 24118 10792 24124 10804
rect 24075 10764 24124 10792
rect 24075 10761 24087 10764
rect 24029 10755 24087 10761
rect 24118 10752 24124 10764
rect 24176 10752 24182 10804
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 6328 10696 6377 10724
rect 6328 10684 6334 10696
rect 6365 10693 6377 10696
rect 6411 10693 6423 10727
rect 6365 10687 6423 10693
rect 19337 10727 19395 10733
rect 19337 10693 19349 10727
rect 19383 10693 19395 10727
rect 19337 10687 19395 10693
rect 21269 10727 21327 10733
rect 21269 10693 21281 10727
rect 21315 10724 21327 10727
rect 21821 10727 21879 10733
rect 21821 10724 21833 10727
rect 21315 10696 21833 10724
rect 21315 10693 21327 10696
rect 21269 10687 21327 10693
rect 21821 10693 21833 10696
rect 21867 10693 21879 10727
rect 21821 10687 21879 10693
rect 24305 10727 24363 10733
rect 24305 10693 24317 10727
rect 24351 10724 24363 10727
rect 25133 10727 25191 10733
rect 25133 10724 25145 10727
rect 24351 10696 25145 10724
rect 24351 10693 24363 10696
rect 24305 10687 24363 10693
rect 25133 10693 25145 10696
rect 25179 10693 25191 10727
rect 25133 10687 25191 10693
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4522 10656 4528 10668
rect 4479 10628 4528 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 8665 10659 8723 10665
rect 4672 10628 6776 10656
rect 4672 10616 4678 10628
rect 5534 10548 5540 10600
rect 5592 10548 5598 10600
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 6748 10529 6776 10628
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8711 10628 8892 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8628 10560 8769 10588
rect 8628 10548 8634 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8864 10588 8892 10628
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9490 10656 9496 10668
rect 9079 10628 9496 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 10928 10628 11529 10656
rect 10928 10616 10934 10628
rect 11517 10625 11529 10628
rect 11563 10656 11575 10659
rect 13541 10659 13599 10665
rect 11563 10628 12434 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 9674 10588 9680 10600
rect 8864 10560 9680 10588
rect 8757 10551 8815 10557
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 12406 10588 12434 10628
rect 13541 10625 13553 10659
rect 13587 10656 13599 10659
rect 13630 10656 13636 10668
rect 13587 10628 13636 10656
rect 13587 10625 13599 10628
rect 13541 10619 13599 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 13817 10659 13875 10665
rect 13817 10656 13829 10659
rect 13771 10628 13829 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 13817 10625 13829 10628
rect 13863 10656 13875 10659
rect 14366 10656 14372 10668
rect 13863 10628 14372 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 14366 10616 14372 10628
rect 14424 10656 14430 10668
rect 14918 10656 14924 10668
rect 14424 10628 14924 10656
rect 14424 10616 14430 10628
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15620 10628 15761 10656
rect 15620 10616 15626 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 18414 10616 18420 10668
rect 18472 10616 18478 10668
rect 18509 10659 18567 10665
rect 18509 10625 18521 10659
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 15286 10588 15292 10600
rect 12406 10560 15292 10588
rect 15286 10548 15292 10560
rect 15344 10588 15350 10600
rect 16298 10588 16304 10600
rect 15344 10560 16304 10588
rect 15344 10548 15350 10560
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 18524 10588 18552 10619
rect 18782 10616 18788 10668
rect 18840 10616 18846 10668
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 18966 10656 18972 10668
rect 18923 10628 18972 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 19058 10616 19064 10668
rect 19116 10656 19122 10668
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 19116 10628 19533 10656
rect 19116 10616 19122 10628
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 18524 10560 19380 10588
rect 6733 10523 6791 10529
rect 5224 10492 6592 10520
rect 5224 10480 5230 10492
rect 2590 10412 2596 10464
rect 2648 10412 2654 10464
rect 2774 10412 2780 10464
rect 2832 10412 2838 10464
rect 4985 10455 5043 10461
rect 4985 10421 4997 10455
rect 5031 10452 5043 10455
rect 5350 10452 5356 10464
rect 5031 10424 5356 10452
rect 5031 10421 5043 10424
rect 4985 10415 5043 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5626 10412 5632 10464
rect 5684 10452 5690 10464
rect 6564 10461 6592 10492
rect 6733 10489 6745 10523
rect 6779 10489 6791 10523
rect 6733 10483 6791 10489
rect 12802 10480 12808 10532
rect 12860 10520 12866 10532
rect 13078 10520 13084 10532
rect 12860 10492 13084 10520
rect 12860 10480 12866 10492
rect 13078 10480 13084 10492
rect 13136 10520 13142 10532
rect 18598 10520 18604 10532
rect 13136 10492 18604 10520
rect 13136 10480 13142 10492
rect 18598 10480 18604 10492
rect 18656 10480 18662 10532
rect 19352 10529 19380 10560
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19628 10588 19656 10619
rect 20990 10616 20996 10668
rect 21048 10656 21054 10668
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 21048 10628 21097 10656
rect 21048 10616 21054 10628
rect 21085 10625 21097 10628
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 21358 10616 21364 10668
rect 21416 10616 21422 10668
rect 21450 10616 21456 10668
rect 21508 10616 21514 10668
rect 22002 10616 22008 10668
rect 22060 10616 22066 10668
rect 22278 10616 22284 10668
rect 22336 10616 22342 10668
rect 23658 10616 23664 10668
rect 23716 10616 23722 10668
rect 23842 10616 23848 10668
rect 23900 10616 23906 10668
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 19484 10560 19656 10588
rect 19484 10548 19490 10560
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 24136 10588 24164 10619
rect 24210 10616 24216 10668
rect 24268 10656 24274 10668
rect 24397 10659 24455 10665
rect 24397 10656 24409 10659
rect 24268 10628 24409 10656
rect 24268 10616 24274 10628
rect 24397 10625 24409 10628
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 24486 10616 24492 10668
rect 24544 10616 24550 10668
rect 24762 10616 24768 10668
rect 24820 10616 24826 10668
rect 24946 10616 24952 10668
rect 25004 10616 25010 10668
rect 24578 10588 24584 10600
rect 23532 10560 24584 10588
rect 23532 10548 23538 10560
rect 24578 10548 24584 10560
rect 24636 10548 24642 10600
rect 19337 10523 19395 10529
rect 19337 10489 19349 10523
rect 19383 10489 19395 10523
rect 19337 10483 19395 10489
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 5684 10424 6193 10452
rect 5684 10412 5690 10424
rect 6181 10421 6193 10424
rect 6227 10421 6239 10455
rect 6181 10415 6239 10421
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 13541 10455 13599 10461
rect 13541 10452 13553 10455
rect 13228 10424 13553 10452
rect 13228 10412 13234 10424
rect 13541 10421 13553 10424
rect 13587 10421 13599 10455
rect 13541 10415 13599 10421
rect 13906 10412 13912 10464
rect 13964 10412 13970 10464
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 15841 10455 15899 10461
rect 15841 10452 15853 10455
rect 15804 10424 15853 10452
rect 15804 10412 15810 10424
rect 15841 10421 15853 10424
rect 15887 10421 15899 10455
rect 15841 10415 15899 10421
rect 18693 10455 18751 10461
rect 18693 10421 18705 10455
rect 18739 10452 18751 10455
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 18739 10424 19257 10452
rect 18739 10421 18751 10424
rect 18693 10415 18751 10421
rect 19245 10421 19257 10424
rect 19291 10452 19303 10455
rect 19702 10452 19708 10464
rect 19291 10424 19708 10452
rect 19291 10421 19303 10424
rect 19245 10415 19303 10421
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 21082 10412 21088 10464
rect 21140 10452 21146 10464
rect 21637 10455 21695 10461
rect 21637 10452 21649 10455
rect 21140 10424 21649 10452
rect 21140 10412 21146 10424
rect 21637 10421 21649 10424
rect 21683 10421 21695 10455
rect 21637 10415 21695 10421
rect 24118 10412 24124 10464
rect 24176 10452 24182 10464
rect 24673 10455 24731 10461
rect 24673 10452 24685 10455
rect 24176 10424 24685 10452
rect 24176 10412 24182 10424
rect 24673 10421 24685 10424
rect 24719 10421 24731 10455
rect 24673 10415 24731 10421
rect 1104 10362 26312 10384
rect 1104 10310 4101 10362
rect 4153 10310 4165 10362
rect 4217 10310 4229 10362
rect 4281 10310 4293 10362
rect 4345 10310 4357 10362
rect 4409 10310 10403 10362
rect 10455 10310 10467 10362
rect 10519 10310 10531 10362
rect 10583 10310 10595 10362
rect 10647 10310 10659 10362
rect 10711 10310 16705 10362
rect 16757 10310 16769 10362
rect 16821 10310 16833 10362
rect 16885 10310 16897 10362
rect 16949 10310 16961 10362
rect 17013 10310 23007 10362
rect 23059 10310 23071 10362
rect 23123 10310 23135 10362
rect 23187 10310 23199 10362
rect 23251 10310 23263 10362
rect 23315 10310 26312 10362
rect 1104 10288 26312 10310
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 6914 10248 6920 10260
rect 6788 10220 6920 10248
rect 6788 10208 6794 10220
rect 6914 10208 6920 10220
rect 6972 10248 6978 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 6972 10220 7297 10248
rect 6972 10208 6978 10220
rect 7285 10217 7297 10220
rect 7331 10217 7343 10251
rect 7285 10211 7343 10217
rect 8938 10208 8944 10260
rect 8996 10248 9002 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8996 10220 9137 10248
rect 8996 10208 9002 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 11974 10208 11980 10260
rect 12032 10208 12038 10260
rect 13538 10208 13544 10260
rect 13596 10248 13602 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 13596 10220 14381 10248
rect 13596 10208 13602 10220
rect 14369 10217 14381 10220
rect 14415 10248 14427 10251
rect 14734 10248 14740 10260
rect 14415 10220 14740 10248
rect 14415 10217 14427 10220
rect 14369 10211 14427 10217
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 15933 10251 15991 10257
rect 15933 10217 15945 10251
rect 15979 10248 15991 10251
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 15979 10220 16405 10248
rect 15979 10217 15991 10220
rect 15933 10211 15991 10217
rect 16393 10217 16405 10220
rect 16439 10248 16451 10251
rect 16942 10248 16948 10260
rect 16439 10220 16948 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 17681 10251 17739 10257
rect 17681 10217 17693 10251
rect 17727 10248 17739 10251
rect 18322 10248 18328 10260
rect 17727 10220 18328 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 18322 10208 18328 10220
rect 18380 10248 18386 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 18380 10220 18429 10248
rect 18380 10208 18386 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 18417 10211 18475 10217
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 19613 10251 19671 10257
rect 19613 10248 19625 10251
rect 18656 10220 19625 10248
rect 18656 10208 18662 10220
rect 19613 10217 19625 10220
rect 19659 10217 19671 10251
rect 20395 10251 20453 10257
rect 20395 10248 20407 10251
rect 19613 10211 19671 10217
rect 20088 10220 20407 10248
rect 2130 10140 2136 10192
rect 2188 10140 2194 10192
rect 13722 10180 13728 10192
rect 12406 10152 13728 10180
rect 2148 10112 2176 10140
rect 2225 10115 2283 10121
rect 2225 10112 2237 10115
rect 2148 10084 2237 10112
rect 2225 10081 2237 10084
rect 2271 10081 2283 10115
rect 12406 10112 12434 10152
rect 13722 10140 13728 10152
rect 13780 10180 13786 10192
rect 15654 10180 15660 10192
rect 13780 10152 15660 10180
rect 13780 10140 13786 10152
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 16853 10183 16911 10189
rect 16853 10149 16865 10183
rect 16899 10180 16911 10183
rect 17034 10180 17040 10192
rect 16899 10152 17040 10180
rect 16899 10149 16911 10152
rect 16853 10143 16911 10149
rect 17034 10140 17040 10152
rect 17092 10180 17098 10192
rect 17313 10183 17371 10189
rect 17313 10180 17325 10183
rect 17092 10152 17325 10180
rect 17092 10140 17098 10152
rect 17313 10149 17325 10152
rect 17359 10149 17371 10183
rect 17313 10143 17371 10149
rect 17865 10183 17923 10189
rect 17865 10149 17877 10183
rect 17911 10180 17923 10183
rect 18506 10180 18512 10192
rect 17911 10152 18512 10180
rect 17911 10149 17923 10152
rect 17865 10143 17923 10149
rect 2225 10075 2283 10081
rect 5276 10084 12434 10112
rect 5276 10056 5304 10084
rect 12802 10072 12808 10124
rect 12860 10072 12866 10124
rect 13354 10112 13360 10124
rect 12912 10084 13360 10112
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10044 2191 10047
rect 2774 10044 2780 10056
rect 2179 10016 2780 10044
rect 2179 10013 2191 10016
rect 2133 10007 2191 10013
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 2470 9979 2528 9985
rect 2470 9976 2482 9979
rect 1964 9948 2482 9976
rect 1964 9917 1992 9948
rect 2470 9945 2482 9948
rect 2516 9945 2528 9979
rect 5000 9976 5028 10007
rect 5166 10004 5172 10056
rect 5224 10004 5230 10056
rect 5258 10004 5264 10056
rect 5316 10004 5322 10056
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 5960 10016 7236 10044
rect 5960 10004 5966 10016
rect 5994 9976 6000 9988
rect 5000 9948 6000 9976
rect 2470 9939 2528 9945
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 6822 9936 6828 9988
rect 6880 9976 6886 9988
rect 7101 9979 7159 9985
rect 7101 9976 7113 9979
rect 6880 9948 7113 9976
rect 6880 9936 6886 9948
rect 7101 9945 7113 9948
rect 7147 9945 7159 9979
rect 7208 9976 7236 10016
rect 7484 10016 7757 10044
rect 7301 9979 7359 9985
rect 7301 9976 7313 9979
rect 7208 9948 7313 9976
rect 7101 9939 7159 9945
rect 7301 9945 7313 9948
rect 7347 9945 7359 9979
rect 7301 9939 7359 9945
rect 1949 9911 2007 9917
rect 1949 9877 1961 9911
rect 1995 9877 2007 9911
rect 1949 9871 2007 9877
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9908 3663 9911
rect 3786 9908 3792 9920
rect 3651 9880 3792 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 6362 9908 6368 9920
rect 5215 9880 6368 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 6546 9868 6552 9920
rect 6604 9868 6610 9920
rect 7484 9917 7512 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 9033 10047 9091 10053
rect 9033 10013 9045 10047
rect 9079 10044 9091 10047
rect 9122 10044 9128 10056
rect 9079 10016 9128 10044
rect 9079 10013 9091 10016
rect 9033 10007 9091 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 9674 10044 9680 10056
rect 9263 10016 9680 10044
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 9674 10004 9680 10016
rect 9732 10044 9738 10056
rect 10962 10044 10968 10056
rect 9732 10016 10968 10044
rect 9732 10004 9738 10016
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10044 11483 10047
rect 11514 10044 11520 10056
rect 11471 10016 11520 10044
rect 11471 10013 11483 10016
rect 11425 10007 11483 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 12526 10004 12532 10056
rect 12584 10004 12590 10056
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 12820 10044 12848 10072
rect 12912 10053 12940 10084
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 13906 10112 13912 10124
rect 13464 10084 13912 10112
rect 12759 10016 12848 10044
rect 12897 10047 12955 10053
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 13170 10004 13176 10056
rect 13228 10004 13234 10056
rect 13464 10053 13492 10084
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 15764 10084 16712 10112
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13688 10016 14289 10044
rect 13688 10004 13694 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14366 10004 14372 10056
rect 14424 10004 14430 10056
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14918 10044 14924 10056
rect 14516 10016 14924 10044
rect 14516 10004 14522 10016
rect 14918 10004 14924 10016
rect 14976 10044 14982 10056
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 14976 10016 15117 10044
rect 14976 10004 14982 10016
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 12860 9948 13308 9976
rect 12860 9936 12866 9948
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9877 7527 9911
rect 7469 9871 7527 9877
rect 7558 9868 7564 9920
rect 7616 9868 7622 9920
rect 12253 9911 12311 9917
rect 12253 9877 12265 9911
rect 12299 9908 12311 9911
rect 13170 9908 13176 9920
rect 12299 9880 13176 9908
rect 12299 9877 12311 9880
rect 12253 9871 12311 9877
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 13280 9908 13308 9948
rect 13354 9936 13360 9988
rect 13412 9936 13418 9988
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 15764 9985 15792 10084
rect 16684 10056 16712 10084
rect 16390 10044 16396 10056
rect 16224 10016 16396 10044
rect 14093 9979 14151 9985
rect 14093 9976 14105 9979
rect 13872 9948 14105 9976
rect 13872 9936 13878 9948
rect 14093 9945 14105 9948
rect 14139 9945 14151 9979
rect 14093 9939 14151 9945
rect 15289 9979 15347 9985
rect 15289 9945 15301 9979
rect 15335 9976 15347 9979
rect 15749 9979 15807 9985
rect 15749 9976 15761 9979
rect 15335 9948 15761 9976
rect 15335 9945 15347 9948
rect 15289 9939 15347 9945
rect 15749 9945 15761 9948
rect 15795 9945 15807 9979
rect 15749 9939 15807 9945
rect 15965 9979 16023 9985
rect 15965 9945 15977 9979
rect 16011 9976 16023 9979
rect 16224 9976 16252 10016
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16666 10004 16672 10056
rect 16724 10004 16730 10056
rect 16011 9948 16252 9976
rect 16011 9945 16023 9948
rect 15965 9939 16023 9945
rect 16298 9936 16304 9988
rect 16356 9936 16362 9988
rect 17328 9976 17356 10143
rect 18506 10140 18512 10152
rect 18564 10140 18570 10192
rect 18432 10084 19196 10112
rect 18432 10053 18460 10084
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10013 18475 10047
rect 18417 10007 18475 10013
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10044 18567 10047
rect 19058 10044 19064 10056
rect 18555 10016 19064 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18138 9976 18144 9988
rect 17328 9948 18144 9976
rect 18138 9936 18144 9948
rect 18196 9976 18202 9988
rect 18524 9976 18552 10007
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 18196 9948 18552 9976
rect 18196 9936 18202 9948
rect 13725 9911 13783 9917
rect 13725 9908 13737 9911
rect 13280 9880 13737 9908
rect 13725 9877 13737 9880
rect 13771 9877 13783 9911
rect 13725 9871 13783 9877
rect 14550 9868 14556 9920
rect 14608 9868 14614 9920
rect 16114 9868 16120 9920
rect 16172 9868 16178 9920
rect 17126 9868 17132 9920
rect 17184 9908 17190 9920
rect 17681 9911 17739 9917
rect 17681 9908 17693 9911
rect 17184 9880 17693 9908
rect 17184 9868 17190 9880
rect 17681 9877 17693 9880
rect 17727 9877 17739 9911
rect 17681 9871 17739 9877
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18104 9880 18797 9908
rect 18104 9868 18110 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 19168 9908 19196 10084
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10044 19303 10047
rect 19702 10044 19708 10056
rect 19291 10016 19708 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 19429 9979 19487 9985
rect 19429 9945 19441 9979
rect 19475 9976 19487 9979
rect 20088 9976 20116 10220
rect 20395 10217 20407 10220
rect 20441 10248 20453 10251
rect 20898 10248 20904 10260
rect 20441 10220 20904 10248
rect 20441 10217 20453 10220
rect 20395 10211 20453 10217
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 22833 10251 22891 10257
rect 22833 10248 22845 10251
rect 21876 10220 22845 10248
rect 21876 10208 21882 10220
rect 22833 10217 22845 10220
rect 22879 10217 22891 10251
rect 22833 10211 22891 10217
rect 20533 10183 20591 10189
rect 20533 10180 20545 10183
rect 19475 9948 20116 9976
rect 20180 10152 20545 10180
rect 19475 9945 19487 9948
rect 19429 9939 19487 9945
rect 20180 9908 20208 10152
rect 20533 10149 20545 10152
rect 20579 10180 20591 10183
rect 20714 10180 20720 10192
rect 20579 10152 20720 10180
rect 20579 10149 20591 10152
rect 20533 10143 20591 10149
rect 20714 10140 20720 10152
rect 20772 10140 20778 10192
rect 20806 10072 20812 10124
rect 20864 10072 20870 10124
rect 21082 10072 21088 10124
rect 21140 10072 21146 10124
rect 22848 10112 22876 10211
rect 22922 10208 22928 10260
rect 22980 10248 22986 10260
rect 23017 10251 23075 10257
rect 23017 10248 23029 10251
rect 22980 10220 23029 10248
rect 22980 10208 22986 10220
rect 23017 10217 23029 10220
rect 23063 10217 23075 10251
rect 23017 10211 23075 10217
rect 24213 10251 24271 10257
rect 24213 10217 24225 10251
rect 24259 10248 24271 10251
rect 24486 10248 24492 10260
rect 24259 10220 24492 10248
rect 24259 10217 24271 10220
rect 24213 10211 24271 10217
rect 24486 10208 24492 10220
rect 24544 10208 24550 10260
rect 24762 10208 24768 10260
rect 24820 10248 24826 10260
rect 24949 10251 25007 10257
rect 24949 10248 24961 10251
rect 24820 10220 24961 10248
rect 24820 10208 24826 10220
rect 24949 10217 24961 10220
rect 24995 10217 25007 10251
rect 24949 10211 25007 10217
rect 23842 10140 23848 10192
rect 23900 10180 23906 10192
rect 25041 10183 25099 10189
rect 25041 10180 25053 10183
rect 23900 10152 25053 10180
rect 23900 10140 23906 10152
rect 23952 10121 23980 10152
rect 25041 10149 25053 10152
rect 25087 10149 25099 10183
rect 25041 10143 25099 10149
rect 23937 10115 23995 10121
rect 22848 10084 23888 10112
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 20272 9976 20300 10007
rect 20622 10004 20628 10056
rect 20680 10044 20686 10056
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 20680 10016 20729 10044
rect 20680 10004 20686 10016
rect 20717 10013 20729 10016
rect 20763 10013 20775 10047
rect 20717 10007 20775 10013
rect 23290 10004 23296 10056
rect 23348 10004 23354 10056
rect 23382 10004 23388 10056
rect 23440 10004 23446 10056
rect 23860 10053 23888 10084
rect 23937 10081 23949 10115
rect 23983 10081 23995 10115
rect 23937 10075 23995 10081
rect 24486 10072 24492 10124
rect 24544 10072 24550 10124
rect 24670 10072 24676 10124
rect 24728 10112 24734 10124
rect 24728 10084 25360 10112
rect 24728 10072 24734 10084
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 24581 10047 24639 10053
rect 23952 10044 24072 10046
rect 24581 10044 24593 10047
rect 23891 10018 24593 10044
rect 23891 10016 23980 10018
rect 24044 10016 24593 10018
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24581 10013 24593 10016
rect 24627 10044 24639 10047
rect 24854 10044 24860 10056
rect 24627 10016 24860 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10044 25099 10047
rect 25130 10044 25136 10056
rect 25087 10016 25136 10044
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25332 10053 25360 10084
rect 25225 10047 25283 10053
rect 25225 10013 25237 10047
rect 25271 10013 25283 10047
rect 25225 10007 25283 10013
rect 25317 10047 25375 10053
rect 25317 10013 25329 10047
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 20990 9976 20996 9988
rect 20272 9948 20996 9976
rect 20990 9936 20996 9948
rect 21048 9936 21054 9988
rect 22370 9976 22376 9988
rect 22310 9948 22376 9976
rect 22370 9936 22376 9948
rect 22428 9936 22434 9988
rect 22649 9979 22707 9985
rect 22649 9945 22661 9979
rect 22695 9945 22707 9979
rect 22649 9939 22707 9945
rect 22865 9979 22923 9985
rect 22865 9945 22877 9979
rect 22911 9976 22923 9979
rect 23569 9979 23627 9985
rect 23569 9976 23581 9979
rect 22911 9948 23581 9976
rect 22911 9945 22923 9948
rect 22865 9939 22923 9945
rect 23569 9945 23581 9948
rect 23615 9976 23627 9979
rect 23658 9976 23664 9988
rect 23615 9948 23664 9976
rect 23615 9945 23627 9948
rect 23569 9939 23627 9945
rect 19168 9880 20208 9908
rect 20717 9911 20775 9917
rect 18785 9871 18843 9877
rect 20717 9877 20729 9911
rect 20763 9908 20775 9911
rect 21358 9908 21364 9920
rect 20763 9880 21364 9908
rect 20763 9877 20775 9880
rect 20717 9871 20775 9877
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 22554 9868 22560 9920
rect 22612 9908 22618 9920
rect 22664 9908 22692 9939
rect 23658 9936 23664 9948
rect 23716 9976 23722 9988
rect 24486 9976 24492 9988
rect 23716 9948 24492 9976
rect 23716 9936 23722 9948
rect 24486 9936 24492 9948
rect 24544 9936 24550 9988
rect 22612 9880 22692 9908
rect 22612 9868 22618 9880
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 25240 9908 25268 10007
rect 23348 9880 25268 9908
rect 23348 9868 23354 9880
rect 25406 9868 25412 9920
rect 25464 9868 25470 9920
rect 1104 9818 26312 9840
rect 1104 9766 4761 9818
rect 4813 9766 4825 9818
rect 4877 9766 4889 9818
rect 4941 9766 4953 9818
rect 5005 9766 5017 9818
rect 5069 9766 11063 9818
rect 11115 9766 11127 9818
rect 11179 9766 11191 9818
rect 11243 9766 11255 9818
rect 11307 9766 11319 9818
rect 11371 9766 17365 9818
rect 17417 9766 17429 9818
rect 17481 9766 17493 9818
rect 17545 9766 17557 9818
rect 17609 9766 17621 9818
rect 17673 9766 23667 9818
rect 23719 9766 23731 9818
rect 23783 9766 23795 9818
rect 23847 9766 23859 9818
rect 23911 9766 23923 9818
rect 23975 9766 26312 9818
rect 1104 9744 26312 9766
rect 6546 9704 6552 9716
rect 2240 9676 6552 9704
rect 1762 9528 1768 9580
rect 1820 9528 1826 9580
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2240 9577 2268 9676
rect 5626 9636 5632 9648
rect 4816 9608 5632 9636
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 2188 9540 2237 9568
rect 2188 9528 2194 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2314 9528 2320 9580
rect 2372 9568 2378 9580
rect 2481 9571 2539 9577
rect 2481 9568 2493 9571
rect 2372 9540 2493 9568
rect 2372 9528 2378 9540
rect 2481 9537 2493 9540
rect 2527 9537 2539 9571
rect 2481 9531 2539 9537
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3844 9540 4077 9568
rect 3844 9528 3850 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 4816 9577 4844 9608
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 5994 9596 6000 9648
rect 6052 9596 6058 9648
rect 6380 9636 6408 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9673 9735 9707
rect 9677 9667 9735 9673
rect 9692 9636 9720 9667
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 14093 9707 14151 9713
rect 14093 9704 14105 9707
rect 13412 9676 14105 9704
rect 13412 9664 13418 9676
rect 14093 9673 14105 9676
rect 14139 9673 14151 9707
rect 16761 9707 16819 9713
rect 16761 9704 16773 9707
rect 14093 9667 14151 9673
rect 16592 9676 16773 9704
rect 6380 9608 8340 9636
rect 9692 9608 11008 9636
rect 4765 9571 4844 9577
rect 4765 9537 4777 9571
rect 4811 9540 4844 9571
rect 4811 9537 4823 9540
rect 4765 9531 4823 9537
rect 4890 9528 4896 9580
rect 4948 9528 4954 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5123 9571 5181 9577
rect 5123 9537 5135 9571
rect 5169 9568 5181 9571
rect 6086 9568 6092 9580
rect 5169 9540 6092 9568
rect 5169 9537 5181 9540
rect 5123 9531 5181 9537
rect 1854 9460 1860 9512
rect 1912 9460 1918 9512
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 5000 9500 5028 9531
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6380 9577 6408 9608
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6632 9571 6690 9577
rect 6632 9537 6644 9571
rect 6678 9568 6690 9571
rect 7558 9568 7564 9580
rect 6678 9540 7564 9568
rect 6678 9537 6690 9540
rect 6632 9531 6690 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8018 9528 8024 9580
rect 8076 9528 8082 9580
rect 8312 9577 8340 9608
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9537 8355 9571
rect 8553 9571 8611 9577
rect 8553 9568 8565 9571
rect 8297 9531 8355 9537
rect 8404 9540 8565 9568
rect 5353 9503 5411 9509
rect 5353 9500 5365 9503
rect 3568 9472 5212 9500
rect 3568 9460 3574 9472
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2498 9364 2504 9376
rect 2087 9336 2504 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3605 9367 3663 9373
rect 3605 9364 3617 9367
rect 3476 9336 3617 9364
rect 3476 9324 3482 9336
rect 3605 9333 3617 9336
rect 3651 9333 3663 9367
rect 3605 9327 3663 9333
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4430 9364 4436 9376
rect 4387 9336 4436 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 5074 9364 5080 9376
rect 4571 9336 5080 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5184 9364 5212 9472
rect 5276 9472 5365 9500
rect 5276 9441 5304 9472
rect 5353 9469 5365 9472
rect 5399 9500 5411 9503
rect 5442 9500 5448 9512
rect 5399 9472 5448 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 8404 9500 8432 9540
rect 8553 9537 8565 9540
rect 8599 9537 8611 9571
rect 8553 9531 8611 9537
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9548 9540 10149 9568
rect 9548 9528 9554 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10870 9568 10876 9580
rect 10275 9540 10876 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 10980 9568 11008 9608
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11756 9608 11989 9636
rect 11756 9596 11762 9608
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 12434 9596 12440 9648
rect 12492 9596 12498 9648
rect 13170 9596 13176 9648
rect 13228 9636 13234 9648
rect 13541 9639 13599 9645
rect 13228 9608 13400 9636
rect 13228 9596 13234 9608
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 10980 9540 11897 9568
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12158 9528 12164 9580
rect 12216 9568 12222 9580
rect 12345 9571 12403 9577
rect 12345 9568 12357 9571
rect 12216 9540 12357 9568
rect 12216 9528 12222 9540
rect 12345 9537 12357 9540
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 13372 9568 13400 9608
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 14461 9639 14519 9645
rect 14461 9636 14473 9639
rect 13587 9608 14473 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 14461 9605 14473 9608
rect 14507 9605 14519 9639
rect 14461 9599 14519 9605
rect 15289 9639 15347 9645
rect 15289 9605 15301 9639
rect 15335 9636 15347 9639
rect 15378 9636 15384 9648
rect 15335 9608 15384 9636
rect 15335 9605 15347 9608
rect 15289 9599 15347 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 15749 9639 15807 9645
rect 15749 9605 15761 9639
rect 15795 9636 15807 9639
rect 16114 9636 16120 9648
rect 15795 9608 16120 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 16114 9596 16120 9608
rect 16172 9596 16178 9648
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13372 9540 13737 9568
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 7852 9472 8432 9500
rect 10413 9503 10471 9509
rect 7852 9441 7880 9472
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 10962 9500 10968 9512
rect 10459 9472 10968 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 10962 9460 10968 9472
rect 11020 9500 11026 9512
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 11020 9472 12081 9500
rect 11020 9460 11026 9472
rect 12069 9469 12081 9472
rect 12115 9500 12127 9503
rect 12544 9500 12572 9528
rect 12115 9472 12572 9500
rect 12115 9469 12127 9472
rect 12069 9463 12127 9469
rect 12802 9460 12808 9512
rect 12860 9500 12866 9512
rect 13924 9500 13952 9531
rect 12860 9472 13952 9500
rect 12860 9460 12866 9472
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9401 5319 9435
rect 5261 9395 5319 9401
rect 7837 9435 7895 9441
rect 7837 9401 7849 9435
rect 7883 9401 7895 9435
rect 7837 9395 7895 9401
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 13449 9435 13507 9441
rect 12952 9404 13400 9432
rect 12952 9392 12958 9404
rect 5810 9364 5816 9376
rect 5184 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 7745 9367 7803 9373
rect 7745 9364 7757 9367
rect 6328 9336 7757 9364
rect 6328 9324 6334 9336
rect 7745 9333 7757 9336
rect 7791 9333 7803 9367
rect 7745 9327 7803 9333
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 10318 9364 10324 9376
rect 9815 9336 10324 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 11517 9367 11575 9373
rect 11517 9333 11529 9367
rect 11563 9364 11575 9367
rect 12342 9364 12348 9376
rect 11563 9336 12348 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 13170 9324 13176 9376
rect 13228 9324 13234 9376
rect 13372 9364 13400 9404
rect 13449 9401 13461 9435
rect 13495 9432 13507 9435
rect 13814 9432 13820 9444
rect 13495 9404 13820 9432
rect 13495 9401 13507 9404
rect 13449 9395 13507 9401
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 14016 9364 14044 9531
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14148 9540 14289 9568
rect 14148 9528 14154 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 14424 9540 14565 9568
rect 14424 9528 14430 9540
rect 14553 9537 14565 9540
rect 14599 9537 14611 9571
rect 14553 9531 14611 9537
rect 14918 9528 14924 9580
rect 14976 9528 14982 9580
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9568 16083 9571
rect 16206 9568 16212 9580
rect 16071 9540 16212 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 16206 9528 16212 9540
rect 16264 9568 16270 9580
rect 16592 9568 16620 9676
rect 16761 9673 16773 9676
rect 16807 9673 16819 9707
rect 18230 9704 18236 9716
rect 16761 9667 16819 9673
rect 17788 9676 18236 9704
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 16724 9608 17141 9636
rect 16724 9596 16730 9608
rect 16776 9577 16804 9608
rect 17129 9605 17141 9608
rect 17175 9605 17187 9639
rect 17129 9599 17187 9605
rect 16264 9540 16620 9568
rect 16761 9571 16819 9577
rect 16264 9528 16270 9540
rect 16761 9537 16773 9571
rect 16807 9537 16819 9571
rect 16761 9531 16819 9537
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 15933 9503 15991 9509
rect 15933 9469 15945 9503
rect 15979 9500 15991 9503
rect 16298 9500 16304 9512
rect 15979 9472 16304 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 16209 9435 16267 9441
rect 16209 9432 16221 9435
rect 14240 9404 16221 9432
rect 14240 9392 14246 9404
rect 16209 9401 16221 9404
rect 16255 9401 16267 9435
rect 16209 9395 16267 9401
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 16868 9432 16896 9531
rect 17144 9500 17172 9599
rect 17218 9596 17224 9648
rect 17276 9636 17282 9648
rect 17788 9645 17816 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 20640 9676 21772 9704
rect 20640 9648 20668 9676
rect 17329 9639 17387 9645
rect 17329 9636 17341 9639
rect 17276 9608 17341 9636
rect 17276 9596 17282 9608
rect 17329 9605 17341 9608
rect 17375 9605 17387 9639
rect 17329 9599 17387 9605
rect 17589 9639 17647 9645
rect 17589 9605 17601 9639
rect 17635 9605 17647 9639
rect 17788 9639 17847 9645
rect 17788 9608 17801 9639
rect 17589 9599 17647 9605
rect 17789 9605 17801 9608
rect 17835 9605 17847 9639
rect 17789 9599 17847 9605
rect 18417 9639 18475 9645
rect 18417 9605 18429 9639
rect 18463 9636 18475 9639
rect 18598 9636 18604 9648
rect 18463 9608 18604 9636
rect 18463 9605 18475 9608
rect 18417 9599 18475 9605
rect 17604 9500 17632 9599
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 18690 9596 18696 9648
rect 18748 9596 18754 9648
rect 19429 9639 19487 9645
rect 19429 9636 19441 9639
rect 18984 9608 19441 9636
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9568 18107 9571
rect 18138 9568 18144 9580
rect 18095 9540 18144 9568
rect 18095 9537 18107 9540
rect 18049 9531 18107 9537
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 18874 9528 18880 9580
rect 18932 9528 18938 9580
rect 18984 9577 19012 9608
rect 19429 9605 19441 9608
rect 19475 9605 19487 9639
rect 19429 9599 19487 9605
rect 20622 9596 20628 9648
rect 20680 9596 20686 9648
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 21744 9636 21772 9676
rect 22094 9664 22100 9716
rect 22152 9704 22158 9716
rect 23382 9704 23388 9716
rect 22152 9676 23388 9704
rect 22152 9664 22158 9676
rect 23382 9664 23388 9676
rect 23440 9664 23446 9716
rect 23845 9639 23903 9645
rect 20772 9608 21680 9636
rect 21744 9608 22324 9636
rect 20772 9596 20778 9608
rect 18969 9571 19027 9577
rect 18969 9537 18981 9571
rect 19015 9537 19027 9571
rect 18969 9531 19027 9537
rect 19150 9528 19156 9580
rect 19208 9528 19214 9580
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 19260 9500 19288 9531
rect 19334 9528 19340 9580
rect 19392 9528 19398 9580
rect 20990 9528 20996 9580
rect 21048 9568 21054 9580
rect 21048 9540 21128 9568
rect 21048 9528 21054 9540
rect 17144 9472 17908 9500
rect 17880 9444 17908 9472
rect 18616 9472 19288 9500
rect 20809 9503 20867 9509
rect 16448 9404 16896 9432
rect 16448 9392 16454 9404
rect 16942 9392 16948 9444
rect 17000 9432 17006 9444
rect 17000 9404 17724 9432
rect 17000 9392 17006 9404
rect 13372 9336 14044 9364
rect 15286 9324 15292 9376
rect 15344 9324 15350 9376
rect 17328 9373 17356 9404
rect 17696 9376 17724 9404
rect 17862 9392 17868 9444
rect 17920 9392 17926 9444
rect 18616 9441 18644 9472
rect 20809 9469 20821 9503
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 18601 9435 18659 9441
rect 18601 9401 18613 9435
rect 18647 9401 18659 9435
rect 18601 9395 18659 9401
rect 18690 9392 18696 9444
rect 18748 9432 18754 9444
rect 20714 9432 20720 9444
rect 18748 9404 20720 9432
rect 18748 9392 18754 9404
rect 20714 9392 20720 9404
rect 20772 9432 20778 9444
rect 20824 9432 20852 9463
rect 20772 9404 20852 9432
rect 21100 9432 21128 9540
rect 21358 9528 21364 9580
rect 21416 9528 21422 9580
rect 21542 9528 21548 9580
rect 21600 9528 21606 9580
rect 21652 9568 21680 9608
rect 21818 9568 21824 9580
rect 21652 9540 21824 9568
rect 21818 9528 21824 9540
rect 21876 9568 21882 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21876 9540 22017 9568
rect 21876 9528 21882 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22094 9528 22100 9580
rect 22152 9528 22158 9580
rect 22296 9577 22324 9608
rect 23845 9605 23857 9639
rect 23891 9636 23903 9639
rect 24118 9636 24124 9648
rect 23891 9608 24124 9636
rect 23891 9605 23903 9608
rect 23845 9599 23903 9605
rect 24118 9596 24124 9608
rect 24176 9596 24182 9648
rect 25406 9636 25412 9648
rect 25070 9608 25412 9636
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9568 22339 9571
rect 22554 9568 22560 9580
rect 22327 9540 22560 9568
rect 22327 9537 22339 9540
rect 22281 9531 22339 9537
rect 22554 9528 22560 9540
rect 22612 9528 22618 9580
rect 21450 9460 21456 9512
rect 21508 9460 21514 9512
rect 22189 9503 22247 9509
rect 22189 9469 22201 9503
rect 22235 9500 22247 9503
rect 22235 9472 22324 9500
rect 22235 9469 22247 9472
rect 22189 9463 22247 9469
rect 22296 9432 22324 9472
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 23569 9503 23627 9509
rect 23569 9500 23581 9503
rect 23440 9472 23581 9500
rect 23440 9460 23446 9472
rect 23569 9469 23581 9472
rect 23615 9469 23627 9503
rect 23569 9463 23627 9469
rect 24854 9460 24860 9512
rect 24912 9500 24918 9512
rect 25593 9503 25651 9509
rect 25593 9500 25605 9503
rect 24912 9472 25605 9500
rect 24912 9460 24918 9472
rect 25593 9469 25605 9472
rect 25639 9469 25651 9503
rect 25593 9463 25651 9469
rect 22462 9432 22468 9444
rect 21100 9404 22468 9432
rect 20772 9392 20778 9404
rect 22462 9392 22468 9404
rect 22520 9432 22526 9444
rect 23290 9432 23296 9444
rect 22520 9404 23296 9432
rect 22520 9392 22526 9404
rect 23290 9392 23296 9404
rect 23348 9392 23354 9444
rect 15473 9367 15531 9373
rect 15473 9333 15485 9367
rect 15519 9364 15531 9367
rect 15749 9367 15807 9373
rect 15749 9364 15761 9367
rect 15519 9336 15761 9364
rect 15519 9333 15531 9336
rect 15473 9327 15531 9333
rect 15749 9333 15761 9336
rect 15795 9333 15807 9367
rect 15749 9327 15807 9333
rect 17313 9367 17371 9373
rect 17313 9333 17325 9367
rect 17359 9333 17371 9367
rect 17313 9327 17371 9333
rect 17494 9324 17500 9376
rect 17552 9324 17558 9376
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17736 9336 17785 9364
rect 17736 9324 17742 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 17957 9367 18015 9373
rect 17957 9333 17969 9367
rect 18003 9364 18015 9367
rect 18322 9364 18328 9376
rect 18003 9336 18328 9364
rect 18003 9333 18015 9336
rect 17957 9327 18015 9333
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 18414 9324 18420 9376
rect 18472 9324 18478 9376
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 19610 9364 19616 9376
rect 18932 9336 19616 9364
rect 18932 9324 18938 9336
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 20990 9324 20996 9376
rect 21048 9324 21054 9376
rect 21177 9367 21235 9373
rect 21177 9333 21189 9367
rect 21223 9364 21235 9367
rect 21542 9364 21548 9376
rect 21223 9336 21548 9364
rect 21223 9333 21235 9336
rect 21177 9327 21235 9333
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 21821 9367 21879 9373
rect 21821 9333 21833 9367
rect 21867 9364 21879 9367
rect 22278 9364 22284 9376
rect 21867 9336 22284 9364
rect 21867 9333 21879 9336
rect 21821 9327 21879 9333
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 25130 9364 25136 9376
rect 23532 9336 25136 9364
rect 23532 9324 23538 9336
rect 25130 9324 25136 9336
rect 25188 9324 25194 9376
rect 1104 9274 26312 9296
rect 1104 9222 4101 9274
rect 4153 9222 4165 9274
rect 4217 9222 4229 9274
rect 4281 9222 4293 9274
rect 4345 9222 4357 9274
rect 4409 9222 10403 9274
rect 10455 9222 10467 9274
rect 10519 9222 10531 9274
rect 10583 9222 10595 9274
rect 10647 9222 10659 9274
rect 10711 9222 16705 9274
rect 16757 9222 16769 9274
rect 16821 9222 16833 9274
rect 16885 9222 16897 9274
rect 16949 9222 16961 9274
rect 17013 9222 23007 9274
rect 23059 9222 23071 9274
rect 23123 9222 23135 9274
rect 23187 9222 23199 9274
rect 23251 9222 23263 9274
rect 23315 9222 26312 9274
rect 1104 9200 26312 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2314 9160 2320 9172
rect 2087 9132 2320 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 2501 9163 2559 9169
rect 2501 9129 2513 9163
rect 2547 9160 2559 9163
rect 2590 9160 2596 9172
rect 2547 9132 2596 9160
rect 2547 9129 2559 9132
rect 2501 9123 2559 9129
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 2866 9120 2872 9172
rect 2924 9120 2930 9172
rect 3510 9160 3516 9172
rect 2976 9132 3516 9160
rect 1762 9052 1768 9104
rect 1820 9092 1826 9104
rect 2976 9092 3004 9132
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 4249 9163 4307 9169
rect 4249 9129 4261 9163
rect 4295 9160 4307 9163
rect 4614 9160 4620 9172
rect 4295 9132 4620 9160
rect 4295 9129 4307 9132
rect 4249 9123 4307 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 6549 9163 6607 9169
rect 6549 9160 6561 9163
rect 4908 9132 6561 9160
rect 1820 9064 3004 9092
rect 1820 9052 1826 9064
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 4430 9092 4436 9104
rect 4212 9064 4436 9092
rect 4212 9052 4218 9064
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 4798 9052 4804 9104
rect 4856 9052 4862 9104
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2682 9024 2688 9036
rect 1912 8996 2688 9024
rect 1912 8984 1918 8996
rect 2682 8984 2688 8996
rect 2740 9024 2746 9036
rect 2740 8996 3372 9024
rect 2740 8984 2746 8996
rect 3344 8965 3372 8996
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 3053 8959 3111 8965
rect 2271 8928 2728 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2314 8848 2320 8900
rect 2372 8848 2378 8900
rect 2498 8848 2504 8900
rect 2556 8897 2562 8900
rect 2556 8891 2575 8897
rect 2563 8857 2575 8891
rect 2556 8851 2575 8857
rect 2556 8848 2562 8851
rect 2700 8829 2728 8928
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 2685 8823 2743 8829
rect 2685 8789 2697 8823
rect 2731 8789 2743 8823
rect 3068 8820 3096 8919
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 4672 8928 4721 8956
rect 4672 8916 4678 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4908 8958 4936 9132
rect 6549 9129 6561 9132
rect 6595 9129 6607 9163
rect 6549 9123 6607 9129
rect 6822 9120 6828 9172
rect 6880 9120 6886 9172
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 8018 9160 8024 9172
rect 7055 9132 8024 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 11241 9163 11299 9169
rect 11241 9129 11253 9163
rect 11287 9160 11299 9163
rect 11514 9160 11520 9172
rect 11287 9132 11520 9160
rect 11287 9129 11299 9132
rect 11241 9123 11299 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 11882 9160 11888 9172
rect 11839 9132 11888 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 12802 9160 12808 9172
rect 12115 9132 12808 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13170 9160 13176 9172
rect 13044 9132 13176 9160
rect 13044 9120 13050 9132
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13320 9132 13553 9160
rect 13320 9120 13326 9132
rect 13541 9129 13553 9132
rect 13587 9160 13599 9163
rect 13998 9160 14004 9172
rect 13587 9132 14004 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14090 9120 14096 9172
rect 14148 9120 14154 9172
rect 14461 9163 14519 9169
rect 14461 9129 14473 9163
rect 14507 9160 14519 9163
rect 16390 9160 16396 9172
rect 14507 9132 16396 9160
rect 14507 9129 14519 9132
rect 14461 9123 14519 9129
rect 5353 9095 5411 9101
rect 5353 9061 5365 9095
rect 5399 9092 5411 9095
rect 5626 9092 5632 9104
rect 5399 9064 5632 9092
rect 5399 9061 5411 9064
rect 5353 9055 5411 9061
rect 5626 9052 5632 9064
rect 5684 9092 5690 9104
rect 11900 9092 11928 9120
rect 13446 9092 13452 9104
rect 5684 9064 6224 9092
rect 11900 9064 12572 9092
rect 5684 9052 5690 9064
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 9024 5135 9027
rect 5902 9024 5908 9036
rect 5123 8996 5908 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 5994 8984 6000 9036
rect 6052 8984 6058 9036
rect 6196 9033 6224 9064
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 8993 6239 9027
rect 6454 9024 6460 9036
rect 6181 8987 6239 8993
rect 6288 8996 6460 9024
rect 4985 8959 5043 8965
rect 4985 8958 4997 8959
rect 4908 8930 4997 8958
rect 4709 8919 4767 8925
rect 4985 8925 4997 8930
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 5704 8964 5762 8965
rect 5704 8959 5724 8964
rect 5704 8956 5716 8959
rect 5307 8928 5672 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8888 3295 8891
rect 3436 8888 3464 8916
rect 3283 8860 3464 8888
rect 3283 8857 3295 8860
rect 3237 8851 3295 8857
rect 3786 8848 3792 8900
rect 3844 8848 3850 8900
rect 3804 8820 3832 8848
rect 3068 8792 3832 8820
rect 2685 8783 2743 8789
rect 5534 8780 5540 8832
rect 5592 8780 5598 8832
rect 5644 8820 5672 8928
rect 5700 8925 5716 8956
rect 5700 8924 5724 8925
rect 5704 8919 5724 8924
rect 5718 8912 5724 8919
rect 5776 8912 5782 8964
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6288 8956 6316 8996
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 8168 8996 9873 9024
rect 8168 8984 8174 8996
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 12434 9024 12440 9036
rect 9861 8987 9919 8993
rect 11072 8996 12440 9024
rect 6135 8928 6316 8956
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 6420 8928 6684 8956
rect 6420 8916 6426 8928
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 6546 8888 6552 8900
rect 6052 8860 6552 8888
rect 6052 8848 6058 8860
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 6656 8897 6684 8928
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 9180 8928 9597 8956
rect 9180 8916 9186 8928
rect 9585 8925 9597 8928
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 11072 8956 11100 8996
rect 12434 8984 12440 8996
rect 12492 8984 12498 9036
rect 9723 8928 11100 8956
rect 11517 8959 11575 8965
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 11517 8925 11529 8959
rect 11563 8956 11575 8959
rect 11698 8956 11704 8968
rect 11563 8928 11704 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 12250 8916 12256 8968
rect 12308 8916 12314 8968
rect 12544 8965 12572 9064
rect 12820 9064 13452 9092
rect 12820 9036 12848 9064
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 14182 9092 14188 9104
rect 13688 9064 14188 9092
rect 13688 9052 13694 9064
rect 14182 9052 14188 9064
rect 14240 9052 14246 9104
rect 12802 8984 12808 9036
rect 12860 8984 12866 9036
rect 13078 9024 13084 9036
rect 12912 8996 13084 9024
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8956 12403 8959
rect 12529 8959 12587 8965
rect 12391 8928 12480 8956
rect 12391 8925 12403 8928
rect 12345 8919 12403 8925
rect 6641 8891 6699 8897
rect 6641 8857 6653 8891
rect 6687 8857 6699 8891
rect 6641 8851 6699 8857
rect 6730 8848 6736 8900
rect 6788 8888 6794 8900
rect 10134 8897 10140 8900
rect 6841 8891 6899 8897
rect 6841 8888 6853 8891
rect 6788 8860 6853 8888
rect 6788 8848 6794 8860
rect 6841 8857 6853 8860
rect 6887 8857 6899 8891
rect 10128 8888 10140 8897
rect 10095 8860 10140 8888
rect 6841 8851 6899 8857
rect 10128 8851 10140 8860
rect 10134 8848 10140 8851
rect 10192 8848 10198 8900
rect 12452 8888 12480 8928
rect 12529 8925 12541 8959
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 12912 8888 12940 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 14476 9024 14504 9123
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 16623 9163 16681 9169
rect 16623 9129 16635 9163
rect 16669 9160 16681 9163
rect 17126 9160 17132 9172
rect 16669 9132 17132 9160
rect 16669 9129 16681 9132
rect 16623 9123 16681 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 18325 9163 18383 9169
rect 18325 9160 18337 9163
rect 17552 9132 18337 9160
rect 17552 9120 17558 9132
rect 18325 9129 18337 9132
rect 18371 9129 18383 9163
rect 18325 9123 18383 9129
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 18601 9163 18659 9169
rect 18601 9160 18613 9163
rect 18472 9132 18613 9160
rect 18472 9120 18478 9132
rect 18601 9129 18613 9132
rect 18647 9160 18659 9163
rect 19334 9160 19340 9172
rect 18647 9132 19340 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 20990 9120 20996 9172
rect 21048 9160 21054 9172
rect 22094 9160 22100 9172
rect 21048 9132 22100 9160
rect 21048 9120 21054 9132
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22281 9163 22339 9169
rect 22281 9129 22293 9163
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 18141 9095 18199 9101
rect 18141 9061 18153 9095
rect 18187 9092 18199 9095
rect 19702 9092 19708 9104
rect 18187 9064 19708 9092
rect 18187 9061 18199 9064
rect 18141 9055 18199 9061
rect 19702 9052 19708 9064
rect 19760 9052 19766 9104
rect 22296 9092 22324 9123
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22557 9163 22615 9169
rect 22557 9160 22569 9163
rect 22428 9132 22569 9160
rect 22428 9120 22434 9132
rect 22557 9129 22569 9132
rect 22603 9129 22615 9163
rect 22557 9123 22615 9129
rect 22462 9092 22468 9104
rect 22296 9064 22468 9092
rect 22462 9052 22468 9064
rect 22520 9052 22526 9104
rect 13320 8996 14504 9024
rect 13320 8984 13326 8996
rect 13372 8965 13400 8996
rect 14826 8984 14832 9036
rect 14884 9024 14890 9036
rect 16574 9024 16580 9036
rect 14884 8996 16580 9024
rect 14884 8984 14890 8996
rect 16574 8984 16580 8996
rect 16632 9024 16638 9036
rect 20533 9027 20591 9033
rect 20533 9024 20545 9027
rect 16632 8996 20545 9024
rect 16632 8984 16638 8996
rect 20533 8993 20545 8996
rect 20579 9024 20591 9027
rect 20806 9024 20812 9036
rect 20579 8996 20812 9024
rect 20579 8993 20591 8996
rect 20533 8987 20591 8993
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 12452 8860 12940 8888
rect 6270 8820 6276 8832
rect 5644 8792 6276 8820
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 11974 8780 11980 8832
rect 12032 8780 12038 8832
rect 13004 8820 13032 8919
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 14056 8928 14289 8956
rect 14056 8916 14062 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 13078 8848 13084 8900
rect 13136 8888 13142 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 13136 8860 13185 8888
rect 13136 8848 13142 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8888 13323 8891
rect 13446 8888 13452 8900
rect 13311 8860 13452 8888
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 13446 8848 13452 8860
rect 13504 8888 13510 8900
rect 14568 8888 14596 8919
rect 15194 8916 15200 8968
rect 15252 8916 15258 8968
rect 18046 8916 18052 8968
rect 18104 8916 18110 8968
rect 18230 8916 18236 8968
rect 18288 8916 18294 8968
rect 18506 8916 18512 8968
rect 18564 8916 18570 8968
rect 18601 8959 18659 8965
rect 18601 8925 18613 8959
rect 18647 8956 18659 8959
rect 18690 8956 18696 8968
rect 18647 8928 18696 8956
rect 18647 8925 18659 8928
rect 18601 8919 18659 8925
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8956 18843 8959
rect 19058 8956 19064 8968
rect 18831 8928 19064 8956
rect 18831 8925 18843 8928
rect 18785 8919 18843 8925
rect 19058 8916 19064 8928
rect 19116 8916 19122 8968
rect 19245 8959 19303 8965
rect 19245 8925 19257 8959
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 13504 8860 14596 8888
rect 13504 8848 13510 8860
rect 15746 8848 15752 8900
rect 15804 8848 15810 8900
rect 17773 8891 17831 8897
rect 17773 8888 17785 8891
rect 16316 8860 17785 8888
rect 13354 8820 13360 8832
rect 13004 8792 13360 8820
rect 13354 8780 13360 8792
rect 13412 8820 13418 8832
rect 16316 8820 16344 8860
rect 17773 8857 17785 8860
rect 17819 8857 17831 8891
rect 18524 8888 18552 8916
rect 19150 8888 19156 8900
rect 18524 8860 19156 8888
rect 17773 8851 17831 8857
rect 19150 8848 19156 8860
rect 19208 8888 19214 8900
rect 19260 8888 19288 8919
rect 19208 8860 19288 8888
rect 19444 8888 19472 8919
rect 20254 8916 20260 8968
rect 20312 8916 20318 8968
rect 22465 8959 22523 8965
rect 22465 8925 22477 8959
rect 22511 8956 22523 8959
rect 22554 8956 22560 8968
rect 22511 8928 22560 8956
rect 22511 8925 22523 8928
rect 22465 8919 22523 8925
rect 22554 8916 22560 8928
rect 22612 8956 22618 8968
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 22612 8928 24409 8956
rect 22612 8916 22618 8928
rect 24397 8925 24409 8928
rect 24443 8956 24455 8959
rect 24670 8956 24676 8968
rect 24443 8928 24676 8956
rect 24443 8925 24455 8928
rect 24397 8919 24455 8925
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 20349 8891 20407 8897
rect 20349 8888 20361 8891
rect 19444 8860 20361 8888
rect 19208 8848 19214 8860
rect 20349 8857 20361 8860
rect 20395 8888 20407 8891
rect 20809 8891 20867 8897
rect 20809 8888 20821 8891
rect 20395 8860 20821 8888
rect 20395 8857 20407 8860
rect 20349 8851 20407 8857
rect 20809 8857 20821 8860
rect 20855 8857 20867 8891
rect 22646 8888 22652 8900
rect 22034 8860 22652 8888
rect 20809 8851 20867 8857
rect 22646 8848 22652 8860
rect 22704 8848 22710 8900
rect 13412 8792 16344 8820
rect 13412 8780 13418 8792
rect 16482 8780 16488 8832
rect 16540 8820 16546 8832
rect 17862 8820 17868 8832
rect 16540 8792 17868 8820
rect 16540 8780 16546 8792
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18138 8780 18144 8832
rect 18196 8820 18202 8832
rect 18969 8823 19027 8829
rect 18969 8820 18981 8823
rect 18196 8792 18981 8820
rect 18196 8780 18202 8792
rect 18969 8789 18981 8792
rect 19015 8789 19027 8823
rect 18969 8783 19027 8789
rect 19334 8780 19340 8832
rect 19392 8780 19398 8832
rect 24394 8780 24400 8832
rect 24452 8820 24458 8832
rect 24489 8823 24547 8829
rect 24489 8820 24501 8823
rect 24452 8792 24501 8820
rect 24452 8780 24458 8792
rect 24489 8789 24501 8792
rect 24535 8789 24547 8823
rect 24489 8783 24547 8789
rect 1104 8730 26312 8752
rect 1104 8678 4761 8730
rect 4813 8678 4825 8730
rect 4877 8678 4889 8730
rect 4941 8678 4953 8730
rect 5005 8678 5017 8730
rect 5069 8678 11063 8730
rect 11115 8678 11127 8730
rect 11179 8678 11191 8730
rect 11243 8678 11255 8730
rect 11307 8678 11319 8730
rect 11371 8678 17365 8730
rect 17417 8678 17429 8730
rect 17481 8678 17493 8730
rect 17545 8678 17557 8730
rect 17609 8678 17621 8730
rect 17673 8678 23667 8730
rect 23719 8678 23731 8730
rect 23783 8678 23795 8730
rect 23847 8678 23859 8730
rect 23911 8678 23923 8730
rect 23975 8678 26312 8730
rect 1104 8656 26312 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1946 8616 1952 8628
rect 1627 8588 1952 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4212 8588 4844 8616
rect 4212 8576 4218 8588
rect 3789 8551 3847 8557
rect 3789 8517 3801 8551
rect 3835 8517 3847 8551
rect 3789 8511 3847 8517
rect 4005 8551 4063 8557
rect 4005 8517 4017 8551
rect 4051 8548 4063 8551
rect 4522 8548 4528 8560
rect 4051 8520 4528 8548
rect 4051 8517 4063 8520
rect 4005 8511 4063 8517
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 3804 8480 3832 8511
rect 4522 8508 4528 8520
rect 4580 8508 4586 8560
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 4709 8551 4767 8557
rect 4709 8548 4721 8551
rect 4672 8520 4721 8548
rect 4672 8508 4678 8520
rect 4709 8517 4721 8520
rect 4755 8517 4767 8551
rect 4816 8548 4844 8588
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 5040 8588 5273 8616
rect 5040 8576 5046 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5442 8616 5448 8628
rect 5261 8579 5319 8585
rect 5368 8588 5448 8616
rect 5368 8548 5396 8588
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 6914 8616 6920 8628
rect 5776 8588 6920 8616
rect 5776 8576 5782 8588
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 9490 8576 9496 8628
rect 9548 8576 9554 8628
rect 12529 8619 12587 8625
rect 12529 8585 12541 8619
rect 12575 8616 12587 8619
rect 13446 8616 13452 8628
rect 12575 8588 13452 8616
rect 12575 8585 12587 8588
rect 12529 8579 12587 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 16298 8576 16304 8628
rect 16356 8576 16362 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 16448 8588 17877 8616
rect 16448 8576 16454 8588
rect 17865 8585 17877 8588
rect 17911 8585 17923 8619
rect 17865 8579 17923 8585
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 20312 8588 22477 8616
rect 20312 8576 20318 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22465 8579 22523 8585
rect 22646 8576 22652 8628
rect 22704 8576 22710 8628
rect 25130 8576 25136 8628
rect 25188 8576 25194 8628
rect 6270 8548 6276 8560
rect 4816 8520 5396 8548
rect 5460 8520 6276 8548
rect 4709 8511 4767 8517
rect 5460 8489 5488 8520
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 11974 8508 11980 8560
rect 12032 8548 12038 8560
rect 12032 8520 12204 8548
rect 12032 8508 12038 8520
rect 5445 8483 5503 8489
rect 3292 8452 4936 8480
rect 3292 8440 3298 8452
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 3252 8412 3280 8440
rect 2372 8384 3280 8412
rect 2372 8372 2378 8384
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 4706 8344 4712 8356
rect 2740 8316 4712 8344
rect 2740 8304 2746 8316
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 3973 8279 4031 8285
rect 3973 8276 3985 8279
rect 2648 8248 3985 8276
rect 2648 8236 2654 8248
rect 3973 8245 3985 8248
rect 4019 8245 4031 8279
rect 3973 8239 4031 8245
rect 4157 8279 4215 8285
rect 4157 8245 4169 8279
rect 4203 8276 4215 8279
rect 4614 8276 4620 8288
rect 4203 8248 4620 8276
rect 4203 8245 4215 8248
rect 4157 8239 4215 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 4908 8276 4936 8452
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8412 5227 8415
rect 5828 8412 5856 8443
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 8386 8489 8392 8492
rect 8380 8443 8392 8489
rect 8386 8440 8392 8443
rect 8444 8440 8450 8492
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 10928 8452 11529 8480
rect 10928 8440 10934 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 12066 8440 12072 8492
rect 12124 8440 12130 8492
rect 12176 8480 12204 8520
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 12802 8548 12808 8560
rect 12492 8520 12808 8548
rect 12492 8508 12498 8520
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 12897 8551 12955 8557
rect 12897 8517 12909 8551
rect 12943 8548 12955 8551
rect 14366 8548 14372 8560
rect 12943 8520 14372 8548
rect 12943 8517 12955 8520
rect 12897 8511 12955 8517
rect 13078 8480 13084 8492
rect 12176 8452 13084 8480
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13354 8480 13360 8492
rect 13219 8452 13360 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 13446 8440 13452 8492
rect 13504 8440 13510 8492
rect 13556 8489 13584 8520
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 16117 8551 16175 8557
rect 16117 8517 16129 8551
rect 16163 8548 16175 8551
rect 16482 8548 16488 8560
rect 16163 8520 16488 8548
rect 16163 8517 16175 8520
rect 16117 8511 16175 8517
rect 16482 8508 16488 8520
rect 16540 8508 16546 8560
rect 16666 8508 16672 8560
rect 16724 8508 16730 8560
rect 18506 8548 18512 8560
rect 16960 8520 18512 8548
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 13906 8440 13912 8492
rect 13964 8440 13970 8492
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15344 8452 15761 8480
rect 15344 8440 15350 8452
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 16960 8489 16988 8520
rect 18506 8508 18512 8520
rect 18564 8548 18570 8560
rect 18564 8520 18644 8548
rect 18564 8508 18570 8520
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16264 8452 16957 8480
rect 16264 8440 16270 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18322 8440 18328 8492
rect 18380 8480 18386 8492
rect 18616 8489 18644 8520
rect 20806 8508 20812 8560
rect 20864 8548 20870 8560
rect 20864 8520 23428 8548
rect 20864 8508 20870 8520
rect 23400 8492 23428 8520
rect 23566 8508 23572 8560
rect 23624 8548 23630 8560
rect 23661 8551 23719 8557
rect 23661 8548 23673 8551
rect 23624 8520 23673 8548
rect 23624 8508 23630 8520
rect 23661 8517 23673 8520
rect 23707 8517 23719 8551
rect 23661 8511 23719 8517
rect 24394 8508 24400 8560
rect 24452 8508 24458 8560
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 18380 8452 18429 8480
rect 18380 8440 18386 8452
rect 18417 8449 18429 8452
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 18840 8452 22094 8480
rect 18840 8440 18846 8452
rect 5215 8384 5856 8412
rect 16761 8415 16819 8421
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 16761 8381 16773 8415
rect 16807 8381 16819 8415
rect 16761 8375 16819 8381
rect 21913 8415 21971 8421
rect 21913 8381 21925 8415
rect 21959 8381 21971 8415
rect 22066 8412 22094 8452
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 23382 8440 23388 8492
rect 23440 8440 23446 8492
rect 25593 8483 25651 8489
rect 25593 8449 25605 8483
rect 25639 8449 25651 8483
rect 25593 8443 25651 8449
rect 25608 8412 25636 8443
rect 22066 8384 25636 8412
rect 21913 8375 21971 8381
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5810 8344 5816 8356
rect 5123 8316 5816 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6822 8344 6828 8356
rect 5920 8316 6828 8344
rect 5920 8276 5948 8316
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 11977 8347 12035 8353
rect 11977 8313 11989 8347
rect 12023 8344 12035 8347
rect 12434 8344 12440 8356
rect 12023 8316 12440 8344
rect 12023 8313 12035 8316
rect 11977 8307 12035 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 14093 8347 14151 8353
rect 14093 8344 14105 8347
rect 12544 8316 14105 8344
rect 4908 8248 5948 8276
rect 11793 8279 11851 8285
rect 11793 8245 11805 8279
rect 11839 8276 11851 8279
rect 11882 8276 11888 8288
rect 11839 8248 11888 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 11882 8236 11888 8248
rect 11940 8276 11946 8288
rect 12161 8279 12219 8285
rect 12161 8276 12173 8279
rect 11940 8248 12173 8276
rect 11940 8236 11946 8248
rect 12161 8245 12173 8248
rect 12207 8245 12219 8279
rect 12161 8239 12219 8245
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12544 8276 12572 8316
rect 14093 8313 14105 8316
rect 14139 8313 14151 8347
rect 16776 8344 16804 8375
rect 18046 8344 18052 8356
rect 16776 8316 18052 8344
rect 14093 8307 14151 8313
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 18233 8347 18291 8353
rect 18233 8313 18245 8347
rect 18279 8344 18291 8347
rect 19150 8344 19156 8356
rect 18279 8316 19156 8344
rect 18279 8313 18291 8316
rect 18233 8307 18291 8313
rect 19150 8304 19156 8316
rect 19208 8304 19214 8356
rect 21928 8344 21956 8375
rect 22462 8344 22468 8356
rect 21928 8316 22468 8344
rect 22462 8304 22468 8316
rect 22520 8304 22526 8356
rect 25866 8304 25872 8356
rect 25924 8304 25930 8356
rect 12308 8248 12572 8276
rect 12308 8236 12314 8248
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 13357 8279 13415 8285
rect 13357 8276 13369 8279
rect 13320 8248 13369 8276
rect 13320 8236 13326 8248
rect 13357 8245 13369 8248
rect 13403 8245 13415 8279
rect 13357 8239 13415 8245
rect 13909 8279 13967 8285
rect 13909 8245 13921 8279
rect 13955 8276 13967 8279
rect 14550 8276 14556 8288
rect 13955 8248 14556 8276
rect 13955 8245 13967 8248
rect 13909 8239 13967 8245
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 16114 8236 16120 8288
rect 16172 8236 16178 8288
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 16669 8279 16727 8285
rect 16669 8276 16681 8279
rect 16264 8248 16681 8276
rect 16264 8236 16270 8248
rect 16669 8245 16681 8248
rect 16715 8245 16727 8279
rect 16669 8239 16727 8245
rect 17126 8236 17132 8288
rect 17184 8236 17190 8288
rect 18322 8236 18328 8288
rect 18380 8236 18386 8288
rect 1104 8186 26312 8208
rect 1104 8134 4101 8186
rect 4153 8134 4165 8186
rect 4217 8134 4229 8186
rect 4281 8134 4293 8186
rect 4345 8134 4357 8186
rect 4409 8134 10403 8186
rect 10455 8134 10467 8186
rect 10519 8134 10531 8186
rect 10583 8134 10595 8186
rect 10647 8134 10659 8186
rect 10711 8134 16705 8186
rect 16757 8134 16769 8186
rect 16821 8134 16833 8186
rect 16885 8134 16897 8186
rect 16949 8134 16961 8186
rect 17013 8134 23007 8186
rect 23059 8134 23071 8186
rect 23123 8134 23135 8186
rect 23187 8134 23199 8186
rect 23251 8134 23263 8186
rect 23315 8134 26312 8186
rect 1104 8112 26312 8134
rect 2590 8032 2596 8084
rect 2648 8072 2654 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 2648 8044 3433 8072
rect 2648 8032 2654 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3421 8035 3479 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5905 8075 5963 8081
rect 4571 8044 5304 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 3099 7976 3801 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 2682 7896 2688 7948
rect 2740 7896 2746 7948
rect 4540 7936 4568 8035
rect 4706 7964 4712 8016
rect 4764 7964 4770 8016
rect 4172 7908 4568 7936
rect 4172 7880 4200 7908
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 3234 7760 3240 7812
rect 3292 7760 3298 7812
rect 3988 7800 4016 7831
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4304 7840 4600 7868
rect 4304 7828 4310 7840
rect 4341 7803 4399 7809
rect 4341 7800 4353 7803
rect 3988 7772 4353 7800
rect 4341 7769 4353 7772
rect 4387 7800 4399 7803
rect 4430 7800 4436 7812
rect 4387 7772 4436 7800
rect 4387 7769 4399 7772
rect 4341 7763 4399 7769
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 4572 7809 4600 7840
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 5276 7877 5304 8044
rect 5905 8041 5917 8075
rect 5951 8041 5963 8075
rect 5905 8035 5963 8041
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 5920 8004 5948 8035
rect 6270 8032 6276 8084
rect 6328 8032 6334 8084
rect 7929 8075 7987 8081
rect 7929 8041 7941 8075
rect 7975 8072 7987 8075
rect 8386 8072 8392 8084
rect 7975 8044 8392 8072
rect 7975 8041 7987 8044
rect 7929 8035 7987 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 10134 8072 10140 8084
rect 9723 8044 10140 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12952 8044 13001 8072
rect 12952 8032 12958 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 6362 8004 6368 8016
rect 5684 7976 6368 8004
rect 5684 7964 5690 7976
rect 6362 7964 6368 7976
rect 6420 7964 6426 8016
rect 10226 8004 10232 8016
rect 9968 7976 10232 8004
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7936 5779 7939
rect 5902 7936 5908 7948
rect 5767 7908 5908 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 5261 7871 5319 7877
rect 5261 7868 5273 7871
rect 5224 7840 5273 7868
rect 5224 7828 5230 7840
rect 5261 7837 5273 7840
rect 5307 7868 5319 7871
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5307 7840 5825 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7708 7840 8125 7868
rect 7708 7828 7714 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9968 7877 9996 7976
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 13740 7936 13768 8035
rect 13906 8032 13912 8084
rect 13964 8032 13970 8084
rect 15381 8075 15439 8081
rect 15381 8041 15393 8075
rect 15427 8072 15439 8075
rect 15470 8072 15476 8084
rect 15427 8044 15476 8072
rect 15427 8041 15439 8044
rect 15381 8035 15439 8041
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 16206 8072 16212 8084
rect 15611 8044 16212 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16632 8044 16957 8072
rect 16632 8032 16638 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 16945 8035 17003 8041
rect 17865 8075 17923 8081
rect 17865 8041 17877 8075
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 15013 8007 15071 8013
rect 15013 7973 15025 8007
rect 15059 8004 15071 8007
rect 16482 8004 16488 8016
rect 15059 7976 16488 8004
rect 15059 7973 15071 7976
rect 15013 7967 15071 7973
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 17880 8004 17908 8035
rect 18046 8032 18052 8084
rect 18104 8032 18110 8084
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18509 8075 18567 8081
rect 18509 8072 18521 8075
rect 18472 8044 18521 8072
rect 18472 8032 18478 8044
rect 18509 8041 18521 8044
rect 18555 8041 18567 8075
rect 18509 8035 18567 8041
rect 19702 8032 19708 8084
rect 19760 8032 19766 8084
rect 18138 8004 18144 8016
rect 17880 7976 18144 8004
rect 18138 7964 18144 7976
rect 18196 7964 18202 8016
rect 18230 7964 18236 8016
rect 18288 8004 18294 8016
rect 18693 8007 18751 8013
rect 18693 8004 18705 8007
rect 18288 7976 18705 8004
rect 18288 7964 18294 7976
rect 18693 7973 18705 7976
rect 18739 7973 18751 8007
rect 18693 7967 18751 7973
rect 19518 7964 19524 8016
rect 19576 7964 19582 8016
rect 19334 7936 19340 7948
rect 10192 7908 10456 7936
rect 10192 7896 10198 7908
rect 10428 7877 10456 7908
rect 13464 7908 19340 7936
rect 9953 7871 10011 7877
rect 9953 7868 9965 7871
rect 9272 7840 9965 7868
rect 9272 7828 9278 7840
rect 9953 7837 9965 7840
rect 9999 7837 10011 7871
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9953 7831 10011 7837
rect 10060 7840 10241 7868
rect 10060 7812 10088 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 13464 7877 13492 7908
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 12492 7840 13185 7868
rect 12492 7828 12498 7840
rect 13173 7837 13185 7840
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7837 13415 7871
rect 13357 7831 13415 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 17126 7868 17132 7880
rect 13449 7831 13507 7837
rect 13556 7840 17132 7868
rect 4557 7803 4615 7809
rect 4557 7769 4569 7803
rect 4603 7800 4615 7803
rect 5074 7800 5080 7812
rect 4603 7772 5080 7800
rect 4603 7769 4615 7772
rect 4557 7763 4615 7769
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 9677 7803 9735 7809
rect 9677 7769 9689 7803
rect 9723 7800 9735 7803
rect 10042 7800 10048 7812
rect 9723 7772 10048 7800
rect 9723 7769 9735 7772
rect 9677 7763 9735 7769
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 11790 7800 11796 7812
rect 10152 7772 11796 7800
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 3437 7735 3495 7741
rect 3437 7732 3449 7735
rect 3191 7704 3449 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 3437 7701 3449 7704
rect 3483 7701 3495 7735
rect 3437 7695 3495 7701
rect 3602 7692 3608 7744
rect 3660 7692 3666 7744
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10152 7732 10180 7772
rect 11790 7760 11796 7772
rect 11848 7760 11854 7812
rect 9916 7704 10180 7732
rect 9916 7692 9922 7704
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 13188 7732 13216 7831
rect 13372 7800 13400 7831
rect 13556 7809 13584 7840
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 17420 7840 17509 7868
rect 13541 7803 13599 7809
rect 13541 7800 13553 7803
rect 13372 7772 13553 7800
rect 13541 7769 13553 7772
rect 13587 7769 13599 7803
rect 13541 7763 13599 7769
rect 15654 7760 15660 7812
rect 15712 7760 15718 7812
rect 17420 7800 17448 7840
rect 17497 7837 17509 7840
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 17920 7840 18153 7868
rect 17920 7828 17926 7840
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 22646 7828 22652 7880
rect 22704 7828 22710 7880
rect 17678 7800 17684 7812
rect 17420 7772 17684 7800
rect 13741 7735 13799 7741
rect 13741 7732 13753 7735
rect 13188 7704 13753 7732
rect 13741 7701 13753 7704
rect 13787 7701 13799 7735
rect 13741 7695 13799 7701
rect 15381 7735 15439 7741
rect 15381 7701 15393 7735
rect 15427 7732 15439 7735
rect 15470 7732 15476 7744
rect 15427 7704 15476 7732
rect 15427 7701 15439 7704
rect 15381 7695 15439 7701
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15562 7692 15568 7744
rect 15620 7732 15626 7744
rect 17420 7732 17448 7772
rect 17678 7760 17684 7772
rect 17736 7800 17742 7812
rect 18414 7800 18420 7812
rect 17736 7772 18420 7800
rect 17736 7760 17742 7772
rect 18414 7760 18420 7772
rect 18472 7800 18478 7812
rect 18966 7800 18972 7812
rect 18472 7772 18972 7800
rect 18472 7760 18478 7772
rect 18966 7760 18972 7772
rect 19024 7800 19030 7812
rect 19245 7803 19303 7809
rect 19245 7800 19257 7803
rect 19024 7772 19257 7800
rect 19024 7760 19030 7772
rect 19245 7769 19257 7772
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 15620 7704 17448 7732
rect 15620 7692 15626 7704
rect 17862 7692 17868 7744
rect 17920 7692 17926 7744
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 18509 7735 18567 7741
rect 18509 7732 18521 7735
rect 18012 7704 18521 7732
rect 18012 7692 18018 7704
rect 18509 7701 18521 7704
rect 18555 7701 18567 7735
rect 18509 7695 18567 7701
rect 21450 7692 21456 7744
rect 21508 7732 21514 7744
rect 23201 7735 23259 7741
rect 23201 7732 23213 7735
rect 21508 7704 23213 7732
rect 21508 7692 21514 7704
rect 23201 7701 23213 7704
rect 23247 7701 23259 7735
rect 23201 7695 23259 7701
rect 1104 7642 26312 7664
rect 1104 7590 4761 7642
rect 4813 7590 4825 7642
rect 4877 7590 4889 7642
rect 4941 7590 4953 7642
rect 5005 7590 5017 7642
rect 5069 7590 11063 7642
rect 11115 7590 11127 7642
rect 11179 7590 11191 7642
rect 11243 7590 11255 7642
rect 11307 7590 11319 7642
rect 11371 7590 17365 7642
rect 17417 7590 17429 7642
rect 17481 7590 17493 7642
rect 17545 7590 17557 7642
rect 17609 7590 17621 7642
rect 17673 7590 23667 7642
rect 23719 7590 23731 7642
rect 23783 7590 23795 7642
rect 23847 7590 23859 7642
rect 23911 7590 23923 7642
rect 23975 7590 26312 7642
rect 1104 7568 26312 7590
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 3973 7531 4031 7537
rect 3973 7497 3985 7531
rect 4019 7528 4031 7531
rect 4430 7528 4436 7540
rect 4019 7500 4436 7528
rect 4019 7497 4031 7500
rect 3973 7491 4031 7497
rect 2332 7460 2360 7491
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 10042 7488 10048 7540
rect 10100 7488 10106 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 11701 7531 11759 7537
rect 11701 7528 11713 7531
rect 10284 7500 11713 7528
rect 10284 7488 10290 7500
rect 11701 7497 11713 7500
rect 11747 7497 11759 7531
rect 11701 7491 11759 7497
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 11848 7500 12081 7528
rect 11848 7488 11854 7500
rect 12069 7497 12081 7500
rect 12115 7497 12127 7531
rect 12069 7491 12127 7497
rect 18322 7488 18328 7540
rect 18380 7528 18386 7540
rect 18601 7531 18659 7537
rect 18601 7528 18613 7531
rect 18380 7500 18613 7528
rect 18380 7488 18386 7500
rect 18601 7497 18613 7500
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 19150 7488 19156 7540
rect 19208 7488 19214 7540
rect 22646 7528 22652 7540
rect 20732 7500 22652 7528
rect 2838 7463 2896 7469
rect 2838 7460 2850 7463
rect 2332 7432 2850 7460
rect 2838 7429 2850 7432
rect 2884 7429 2896 7463
rect 2838 7423 2896 7429
rect 10134 7420 10140 7472
rect 10192 7460 10198 7472
rect 10873 7463 10931 7469
rect 10873 7460 10885 7463
rect 10192 7432 10885 7460
rect 10192 7420 10198 7432
rect 10873 7429 10885 7432
rect 10919 7429 10931 7463
rect 11073 7463 11131 7469
rect 11073 7460 11085 7463
rect 10873 7423 10931 7429
rect 10980 7432 11085 7460
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3602 7392 3608 7404
rect 2547 7364 3608 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4212 7364 4261 7392
rect 4212 7352 4218 7364
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 4893 7395 4951 7401
rect 4893 7392 4905 7395
rect 4672 7364 4905 7392
rect 4672 7352 4678 7364
rect 4893 7361 4905 7364
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8168 7364 8217 7392
rect 8168 7352 8174 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8472 7395 8530 7401
rect 8472 7361 8484 7395
rect 8518 7392 8530 7395
rect 8938 7392 8944 7404
rect 8518 7364 8944 7392
rect 8518 7361 8530 7364
rect 8472 7355 8530 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10781 7395 10839 7401
rect 10781 7392 10793 7395
rect 9907 7364 10793 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10781 7361 10793 7364
rect 10827 7392 10839 7395
rect 10980 7392 11008 7432
rect 11073 7429 11085 7432
rect 11119 7429 11131 7463
rect 12250 7460 12256 7472
rect 11073 7423 11131 7429
rect 11532 7432 12256 7460
rect 11532 7401 11560 7432
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 15286 7420 15292 7472
rect 15344 7460 15350 7472
rect 16298 7460 16304 7472
rect 15344 7432 16304 7460
rect 15344 7420 15350 7432
rect 16298 7420 16304 7432
rect 16356 7460 16362 7472
rect 18414 7460 18420 7472
rect 16356 7432 18420 7460
rect 16356 7420 16362 7432
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 18506 7420 18512 7472
rect 18564 7460 18570 7472
rect 18693 7463 18751 7469
rect 18693 7460 18705 7463
rect 18564 7432 18705 7460
rect 18564 7420 18570 7432
rect 18693 7429 18705 7432
rect 18739 7429 18751 7463
rect 18693 7423 18751 7429
rect 19794 7420 19800 7472
rect 19852 7460 19858 7472
rect 20732 7460 20760 7500
rect 22646 7488 22652 7500
rect 22704 7528 22710 7540
rect 23615 7531 23673 7537
rect 23615 7528 23627 7531
rect 22704 7500 23627 7528
rect 22704 7488 22710 7500
rect 23615 7497 23627 7500
rect 23661 7497 23673 7531
rect 23615 7491 23673 7497
rect 19852 7432 20760 7460
rect 19852 7420 19858 7432
rect 10827 7364 11008 7392
rect 11517 7395 11575 7401
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 11517 7361 11529 7395
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 2608 7188 2636 7287
rect 4338 7284 4344 7336
rect 4396 7284 4402 7336
rect 9784 7268 9812 7355
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 12434 7392 12440 7404
rect 11940 7364 12440 7392
rect 11940 7352 11946 7364
rect 12434 7352 12440 7364
rect 12492 7392 12498 7404
rect 12710 7392 12716 7404
rect 12492 7364 12716 7392
rect 12492 7352 12498 7364
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 20732 7401 20760 7432
rect 22554 7420 22560 7472
rect 22612 7420 22618 7472
rect 24026 7420 24032 7472
rect 24084 7460 24090 7472
rect 24670 7460 24676 7472
rect 24084 7432 24676 7460
rect 24084 7420 24090 7432
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 17920 7364 18061 7392
rect 17920 7352 17926 7364
rect 18049 7361 18061 7364
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 21910 7392 21916 7404
rect 21867 7364 21916 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 23753 7395 23811 7401
rect 23753 7361 23765 7395
rect 23799 7392 23811 7395
rect 24302 7392 24308 7404
rect 23799 7364 24308 7392
rect 23799 7361 23811 7364
rect 23753 7355 23811 7361
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 10226 7284 10232 7336
rect 10284 7284 10290 7336
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19518 7324 19524 7336
rect 19392 7296 19524 7324
rect 19392 7284 19398 7296
rect 19518 7284 19524 7296
rect 19576 7324 19582 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 19576 7296 20545 7324
rect 19576 7284 19582 7296
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 20622 7284 20628 7336
rect 20680 7284 20686 7336
rect 20806 7284 20812 7336
rect 20864 7284 20870 7336
rect 21545 7327 21603 7333
rect 21545 7293 21557 7327
rect 21591 7324 21603 7327
rect 22189 7327 22247 7333
rect 22189 7324 22201 7327
rect 21591 7296 22201 7324
rect 21591 7293 21603 7296
rect 21545 7287 21603 7293
rect 22189 7293 22201 7296
rect 22235 7293 22247 7327
rect 22189 7287 22247 7293
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 4617 7259 4675 7265
rect 4617 7256 4629 7259
rect 4580 7228 4629 7256
rect 4580 7216 4586 7228
rect 4617 7225 4629 7228
rect 4663 7225 4675 7259
rect 4617 7219 4675 7225
rect 9766 7216 9772 7268
rect 9824 7256 9830 7268
rect 9824 7228 11100 7256
rect 9824 7216 9830 7228
rect 3786 7188 3792 7200
rect 2608 7160 3792 7188
rect 3786 7148 3792 7160
rect 3844 7148 3850 7200
rect 4706 7148 4712 7200
rect 4764 7148 4770 7200
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 9214 7188 9220 7200
rect 7524 7160 9220 7188
rect 7524 7148 7530 7160
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9582 7148 9588 7200
rect 9640 7148 9646 7200
rect 11072 7197 11100 7228
rect 19058 7216 19064 7268
rect 19116 7216 19122 7268
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 11204 7160 11253 7188
rect 11204 7148 11210 7160
rect 11241 7157 11253 7160
rect 11287 7188 11299 7191
rect 11514 7188 11520 7200
rect 11287 7160 11520 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 17954 7188 17960 7200
rect 16172 7160 17960 7188
rect 16172 7148 16178 7160
rect 17954 7148 17960 7160
rect 18012 7188 18018 7200
rect 18230 7188 18236 7200
rect 18012 7160 18236 7188
rect 18012 7148 18018 7160
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 18417 7191 18475 7197
rect 18417 7157 18429 7191
rect 18463 7188 18475 7191
rect 18506 7188 18512 7200
rect 18463 7160 18512 7188
rect 18463 7157 18475 7160
rect 18417 7151 18475 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 20349 7191 20407 7197
rect 20349 7157 20361 7191
rect 20395 7188 20407 7191
rect 21266 7188 21272 7200
rect 20395 7160 21272 7188
rect 20395 7157 20407 7160
rect 20349 7151 20407 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 1104 7098 26312 7120
rect 1104 7046 4101 7098
rect 4153 7046 4165 7098
rect 4217 7046 4229 7098
rect 4281 7046 4293 7098
rect 4345 7046 4357 7098
rect 4409 7046 10403 7098
rect 10455 7046 10467 7098
rect 10519 7046 10531 7098
rect 10583 7046 10595 7098
rect 10647 7046 10659 7098
rect 10711 7046 16705 7098
rect 16757 7046 16769 7098
rect 16821 7046 16833 7098
rect 16885 7046 16897 7098
rect 16949 7046 16961 7098
rect 17013 7046 23007 7098
rect 23059 7046 23071 7098
rect 23123 7046 23135 7098
rect 23187 7046 23199 7098
rect 23251 7046 23263 7098
rect 23315 7046 26312 7098
rect 1104 7024 26312 7046
rect 5166 6944 5172 6996
rect 5224 6944 5230 6996
rect 5442 6944 5448 6996
rect 5500 6984 5506 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 5500 6956 6101 6984
rect 5500 6944 5506 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 6104 6916 6132 6947
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 6420 6956 6469 6984
rect 6420 6944 6426 6956
rect 6457 6953 6469 6956
rect 6503 6984 6515 6987
rect 7374 6984 7380 6996
rect 6503 6956 7380 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 7466 6944 7472 6996
rect 7524 6944 7530 6996
rect 7650 6944 7656 6996
rect 7708 6944 7714 6996
rect 9125 6987 9183 6993
rect 9125 6984 9137 6987
rect 8680 6956 9137 6984
rect 8680 6925 8708 6956
rect 9125 6953 9137 6956
rect 9171 6953 9183 6987
rect 9125 6947 9183 6953
rect 9493 6987 9551 6993
rect 9493 6953 9505 6987
rect 9539 6984 9551 6987
rect 9766 6984 9772 6996
rect 9539 6956 9772 6984
rect 9539 6953 9551 6956
rect 9493 6947 9551 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 10781 6987 10839 6993
rect 10781 6953 10793 6987
rect 10827 6984 10839 6987
rect 10962 6984 10968 6996
rect 10827 6956 10968 6984
rect 10827 6953 10839 6956
rect 10781 6947 10839 6953
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 12250 6984 12256 6996
rect 11072 6956 12256 6984
rect 8665 6919 8723 6925
rect 8665 6916 8677 6919
rect 6104 6888 8677 6916
rect 8665 6885 8677 6888
rect 8711 6885 8723 6919
rect 8665 6879 8723 6885
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 7006 6848 7012 6860
rect 6319 6820 7012 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 9582 6808 9588 6860
rect 9640 6808 9646 6860
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10873 6851 10931 6857
rect 10873 6848 10885 6851
rect 10376 6820 10885 6848
rect 10376 6808 10382 6820
rect 10873 6817 10885 6820
rect 10919 6817 10931 6851
rect 11072 6848 11100 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 15102 6944 15108 6996
rect 15160 6993 15166 6996
rect 15160 6987 15209 6993
rect 15160 6953 15163 6987
rect 15197 6984 15209 6987
rect 15378 6984 15384 6996
rect 15197 6956 15384 6984
rect 15197 6953 15209 6956
rect 15160 6947 15209 6953
rect 15160 6944 15166 6947
rect 15378 6944 15384 6956
rect 15436 6984 15442 6996
rect 15838 6984 15844 6996
rect 15436 6956 15844 6984
rect 15436 6944 15442 6956
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 16206 6944 16212 6996
rect 16264 6984 16270 6996
rect 18279 6987 18337 6993
rect 16264 6956 18092 6984
rect 16264 6944 16270 6956
rect 15289 6919 15347 6925
rect 15289 6885 15301 6919
rect 15335 6916 15347 6919
rect 16114 6916 16120 6928
rect 15335 6888 16120 6916
rect 15335 6885 15347 6888
rect 15289 6879 15347 6885
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 18064 6916 18092 6956
rect 18279 6953 18291 6987
rect 18325 6984 18337 6987
rect 18414 6984 18420 6996
rect 18325 6956 18420 6984
rect 18325 6953 18337 6956
rect 18279 6947 18337 6953
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 18877 6987 18935 6993
rect 18877 6953 18889 6987
rect 18923 6984 18935 6987
rect 19242 6984 19248 6996
rect 18923 6956 19248 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 20530 6984 20536 6996
rect 19352 6956 20536 6984
rect 18739 6919 18797 6925
rect 18739 6916 18751 6919
rect 18064 6888 18751 6916
rect 18739 6885 18751 6888
rect 18785 6916 18797 6919
rect 19352 6916 19380 6956
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 20806 6944 20812 6996
rect 20864 6984 20870 6996
rect 21131 6987 21189 6993
rect 21131 6984 21143 6987
rect 20864 6956 21143 6984
rect 20864 6944 20870 6956
rect 21131 6953 21143 6956
rect 21177 6953 21189 6987
rect 21131 6947 21189 6953
rect 18785 6888 19380 6916
rect 18785 6885 18797 6888
rect 18739 6879 18797 6885
rect 10873 6811 10931 6817
rect 10980 6820 11100 6848
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5592 6752 5825 6780
rect 5592 6740 5598 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 7098 6780 7104 6792
rect 6963 6752 7104 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 4056 6715 4114 6721
rect 4056 6681 4068 6715
rect 4102 6712 4114 6715
rect 4706 6712 4712 6724
rect 4102 6684 4712 6712
rect 4102 6681 4114 6684
rect 4056 6675 4114 6681
rect 4706 6672 4712 6684
rect 4764 6672 4770 6724
rect 6380 6712 6408 6743
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8343 6752 9045 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 9033 6749 9045 6752
rect 9079 6780 9091 6783
rect 9600 6780 9628 6808
rect 10980 6780 11008 6820
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 12952 6820 16497 6848
rect 12952 6808 12958 6820
rect 16485 6817 16497 6820
rect 16531 6848 16543 6851
rect 17770 6848 17776 6860
rect 16531 6820 17776 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 17770 6808 17776 6820
rect 17828 6848 17834 6860
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 17828 6820 19349 6848
rect 17828 6808 17834 6820
rect 19337 6817 19349 6820
rect 19383 6848 19395 6851
rect 21910 6848 21916 6860
rect 19383 6820 21916 6848
rect 19383 6817 19395 6820
rect 19337 6811 19395 6817
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 22373 6851 22431 6857
rect 22373 6817 22385 6851
rect 22419 6848 22431 6851
rect 22554 6848 22560 6860
rect 22419 6820 22560 6848
rect 22419 6817 22431 6820
rect 22373 6811 22431 6817
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 9079 6752 9628 6780
rect 10888 6752 11008 6780
rect 11057 6783 11115 6789
rect 9079 6749 9091 6752
rect 9033 6743 9091 6749
rect 7190 6712 7196 6724
rect 6380 6684 7196 6712
rect 7190 6672 7196 6684
rect 7248 6672 7254 6724
rect 7285 6715 7343 6721
rect 7285 6681 7297 6715
rect 7331 6712 7343 6715
rect 9306 6712 9312 6724
rect 7331 6684 9312 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 9306 6672 9312 6684
rect 9364 6672 9370 6724
rect 10505 6715 10563 6721
rect 10505 6681 10517 6715
rect 10551 6712 10563 6715
rect 10888 6712 10916 6752
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 12621 6783 12679 6789
rect 11103 6752 12434 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 10551 6684 10916 6712
rect 10551 6681 10563 6684
rect 10505 6675 10563 6681
rect 10962 6672 10968 6724
rect 11020 6672 11026 6724
rect 11324 6715 11382 6721
rect 11324 6681 11336 6715
rect 11370 6712 11382 6715
rect 12158 6712 12164 6724
rect 11370 6684 12164 6712
rect 11370 6681 11382 6684
rect 11324 6675 11382 6681
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 12406 6712 12434 6752
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 12710 6780 12716 6792
rect 12667 6752 12716 6780
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 12894 6712 12900 6724
rect 12406 6684 12900 6712
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 13648 6712 13676 6743
rect 14366 6740 14372 6792
rect 14424 6780 14430 6792
rect 15013 6783 15071 6789
rect 15013 6780 15025 6783
rect 14424 6752 15025 6780
rect 14424 6740 14430 6752
rect 15013 6749 15025 6752
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 14921 6715 14979 6721
rect 14921 6712 14933 6715
rect 13648 6684 14933 6712
rect 14921 6681 14933 6684
rect 14967 6681 14979 6715
rect 15028 6712 15056 6743
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15473 6783 15531 6789
rect 15473 6780 15485 6783
rect 15344 6752 15485 6780
rect 15344 6740 15350 6752
rect 15473 6749 15485 6752
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6780 15715 6783
rect 15746 6780 15752 6792
rect 15703 6752 15752 6780
rect 15703 6749 15715 6752
rect 15657 6743 15715 6749
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 16022 6740 16028 6792
rect 16080 6740 16086 6792
rect 16853 6783 16911 6789
rect 16853 6780 16865 6783
rect 16592 6752 16865 6780
rect 15028 6684 15516 6712
rect 14921 6675 14979 6681
rect 15488 6656 15516 6684
rect 15562 6672 15568 6724
rect 15620 6712 15626 6724
rect 15841 6715 15899 6721
rect 15841 6712 15853 6715
rect 15620 6684 15853 6712
rect 15620 6672 15626 6684
rect 15841 6681 15853 6684
rect 15887 6681 15899 6715
rect 15841 6675 15899 6681
rect 15933 6715 15991 6721
rect 15933 6681 15945 6715
rect 15979 6712 15991 6715
rect 16482 6712 16488 6724
rect 15979 6684 16488 6712
rect 15979 6681 15991 6684
rect 15933 6675 15991 6681
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 6546 6604 6552 6656
rect 6604 6644 6610 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6604 6616 6837 6644
rect 6604 6604 6610 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7009 6647 7067 6653
rect 7009 6644 7021 6647
rect 6972 6616 7021 6644
rect 6972 6604 6978 6616
rect 7009 6613 7021 6616
rect 7055 6613 7067 6647
rect 7009 6607 7067 6613
rect 7495 6647 7553 6653
rect 7495 6613 7507 6647
rect 7541 6644 7553 6647
rect 7834 6644 7840 6656
rect 7541 6616 7840 6644
rect 7541 6613 7553 6616
rect 7495 6607 7553 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9398 6644 9404 6656
rect 8803 6616 9404 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 9732 6616 10241 6644
rect 9732 6604 9738 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10229 6607 10287 6613
rect 10597 6647 10655 6653
rect 10597 6613 10609 6647
rect 10643 6644 10655 6647
rect 11882 6644 11888 6656
rect 10643 6616 11888 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12032 6616 12449 6644
rect 12032 6604 12038 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 13170 6604 13176 6656
rect 13228 6604 13234 6656
rect 13262 6604 13268 6656
rect 13320 6644 13326 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13320 6616 13737 6644
rect 13320 6604 13326 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 15381 6647 15439 6653
rect 15381 6644 15393 6647
rect 15068 6616 15393 6644
rect 15068 6604 15074 6616
rect 15381 6613 15393 6616
rect 15427 6613 15439 6647
rect 15381 6607 15439 6613
rect 15470 6604 15476 6656
rect 15528 6604 15534 6656
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16592 6644 16620 6752
rect 16853 6749 16865 6752
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 18138 6740 18144 6792
rect 18196 6780 18202 6792
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18196 6752 18613 6780
rect 18196 6740 18202 6752
rect 18601 6749 18613 6752
rect 18647 6749 18659 6783
rect 18601 6743 18659 6749
rect 17862 6672 17868 6724
rect 17920 6672 17926 6724
rect 18616 6712 18644 6743
rect 19058 6740 19064 6792
rect 19116 6740 19122 6792
rect 19702 6740 19708 6792
rect 19760 6740 19766 6792
rect 21174 6740 21180 6792
rect 21232 6780 21238 6792
rect 21269 6783 21327 6789
rect 21269 6780 21281 6783
rect 21232 6752 21281 6780
rect 21232 6740 21238 6752
rect 21269 6749 21281 6752
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 22281 6783 22339 6789
rect 22281 6749 22293 6783
rect 22327 6780 22339 6783
rect 23753 6783 23811 6789
rect 23753 6780 23765 6783
rect 22327 6752 23765 6780
rect 22327 6749 22339 6752
rect 22281 6743 22339 6749
rect 23753 6749 23765 6752
rect 23799 6780 23811 6783
rect 24026 6780 24032 6792
rect 23799 6752 24032 6780
rect 23799 6749 23811 6752
rect 23753 6743 23811 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 21361 6715 21419 6721
rect 21361 6712 21373 6715
rect 18616 6684 19380 6712
rect 20746 6684 21373 6712
rect 16255 6616 16620 6644
rect 19061 6647 19119 6653
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 19061 6613 19073 6647
rect 19107 6644 19119 6647
rect 19242 6644 19248 6656
rect 19107 6616 19248 6644
rect 19107 6613 19119 6616
rect 19061 6607 19119 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19352 6644 19380 6684
rect 21361 6681 21373 6684
rect 21407 6681 21419 6715
rect 21361 6675 21419 6681
rect 19794 6644 19800 6656
rect 19352 6616 19800 6644
rect 19794 6604 19800 6616
rect 19852 6604 19858 6656
rect 23566 6604 23572 6656
rect 23624 6644 23630 6656
rect 23845 6647 23903 6653
rect 23845 6644 23857 6647
rect 23624 6616 23857 6644
rect 23624 6604 23630 6616
rect 23845 6613 23857 6616
rect 23891 6613 23903 6647
rect 23845 6607 23903 6613
rect 24118 6604 24124 6656
rect 24176 6604 24182 6656
rect 1104 6554 26312 6576
rect 1104 6502 4761 6554
rect 4813 6502 4825 6554
rect 4877 6502 4889 6554
rect 4941 6502 4953 6554
rect 5005 6502 5017 6554
rect 5069 6502 11063 6554
rect 11115 6502 11127 6554
rect 11179 6502 11191 6554
rect 11243 6502 11255 6554
rect 11307 6502 11319 6554
rect 11371 6502 17365 6554
rect 17417 6502 17429 6554
rect 17481 6502 17493 6554
rect 17545 6502 17557 6554
rect 17609 6502 17621 6554
rect 17673 6502 23667 6554
rect 23719 6502 23731 6554
rect 23783 6502 23795 6554
rect 23847 6502 23859 6554
rect 23911 6502 23923 6554
rect 23975 6502 26312 6554
rect 1104 6480 26312 6502
rect 5534 6440 5540 6452
rect 5000 6412 5540 6440
rect 5000 6381 5028 6412
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5828 6412 6377 6440
rect 5828 6381 5856 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6638 6400 6644 6452
rect 6696 6400 6702 6452
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 6880 6412 7788 6440
rect 6880 6400 6886 6412
rect 4985 6375 5043 6381
rect 4985 6341 4997 6375
rect 5031 6341 5043 6375
rect 4985 6335 5043 6341
rect 5813 6375 5871 6381
rect 5813 6341 5825 6375
rect 5859 6341 5871 6375
rect 5813 6335 5871 6341
rect 5905 6375 5963 6381
rect 5905 6341 5917 6375
rect 5951 6372 5963 6375
rect 6656 6372 6684 6400
rect 5951 6344 6684 6372
rect 6733 6375 6791 6381
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 6733 6341 6745 6375
rect 6779 6372 6791 6375
rect 7650 6372 7656 6384
rect 6779 6344 7656 6372
rect 6779 6341 6791 6344
rect 6733 6335 6791 6341
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 5718 6313 5724 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5685 6307 5724 6313
rect 5685 6273 5697 6307
rect 5685 6267 5724 6273
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5552 6236 5580 6267
rect 5718 6264 5724 6267
rect 5776 6264 5782 6316
rect 6086 6313 6092 6316
rect 6043 6307 6092 6313
rect 6043 6273 6055 6307
rect 6089 6273 6092 6307
rect 6043 6267 6092 6273
rect 6086 6264 6092 6267
rect 6144 6264 6150 6316
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 6822 6304 6828 6316
rect 6687 6276 6828 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6656 6236 6684 6267
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7055 6276 7604 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 5491 6208 5580 6236
rect 5644 6208 6684 6236
rect 6932 6236 6960 6267
rect 7101 6239 7159 6245
rect 6932 6208 7052 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5644 6180 5672 6208
rect 5350 6128 5356 6180
rect 5408 6128 5414 6180
rect 5626 6128 5632 6180
rect 5684 6128 5690 6180
rect 6178 6128 6184 6180
rect 6236 6128 6242 6180
rect 7024 6100 7052 6208
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7282 6236 7288 6248
rect 7147 6208 7288 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7576 6245 7604 6276
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6205 7619 6239
rect 7760 6236 7788 6412
rect 8938 6400 8944 6452
rect 8996 6400 9002 6452
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9214 6440 9220 6452
rect 9171 6412 9220 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9858 6440 9864 6452
rect 9364 6412 9864 6440
rect 9364 6400 9370 6412
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10134 6400 10140 6452
rect 10192 6400 10198 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 10284 6412 10333 6440
rect 10284 6400 10290 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 11974 6440 11980 6452
rect 10321 6403 10379 6409
rect 10796 6412 11980 6440
rect 8389 6375 8447 6381
rect 8389 6341 8401 6375
rect 8435 6372 8447 6375
rect 10152 6372 10180 6400
rect 10796 6372 10824 6412
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12158 6400 12164 6452
rect 12216 6400 12222 6452
rect 15105 6443 15163 6449
rect 15105 6409 15117 6443
rect 15151 6440 15163 6443
rect 15930 6440 15936 6452
rect 15151 6412 15936 6440
rect 15151 6409 15163 6412
rect 15105 6403 15163 6409
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16114 6440 16120 6452
rect 16040 6412 16120 6440
rect 11333 6375 11391 6381
rect 11333 6372 11345 6375
rect 8435 6344 10824 6372
rect 10888 6344 11345 6372
rect 8435 6341 8447 6344
rect 8389 6335 8447 6341
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 8294 6304 8300 6316
rect 7883 6276 8300 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 9122 6307 9180 6313
rect 9122 6273 9134 6307
rect 9168 6304 9180 6307
rect 9306 6304 9312 6316
rect 9168 6276 9312 6304
rect 9168 6273 9180 6276
rect 9122 6267 9180 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9456 6276 9689 6304
rect 9456 6264 9462 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 9825 6307 9883 6313
rect 9825 6273 9837 6307
rect 9871 6304 9883 6307
rect 9871 6273 9904 6304
rect 9825 6267 9904 6273
rect 9585 6239 9643 6245
rect 7760 6208 8708 6236
rect 7561 6199 7619 6205
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 8570 6168 8576 6180
rect 7432 6140 8576 6168
rect 7432 6128 7438 6140
rect 7558 6100 7564 6112
rect 7024 6072 7564 6100
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7944 6109 7972 6140
rect 8570 6128 8576 6140
rect 8628 6128 8634 6180
rect 8680 6177 8708 6208
rect 9585 6205 9597 6239
rect 9631 6236 9643 6239
rect 9631 6208 9812 6236
rect 9631 6205 9643 6208
rect 9585 6199 9643 6205
rect 8665 6171 8723 6177
rect 8665 6137 8677 6171
rect 8711 6137 8723 6171
rect 8665 6131 8723 6137
rect 9493 6171 9551 6177
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 9674 6168 9680 6180
rect 9539 6140 9680 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6069 7987 6103
rect 7929 6063 7987 6069
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 8754 6100 8760 6112
rect 8343 6072 8760 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 8846 6060 8852 6112
rect 8904 6060 8910 6112
rect 9784 6100 9812 6208
rect 9876 6168 9904 6267
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 10226 6313 10232 6316
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10183 6307 10232 6313
rect 10183 6273 10195 6307
rect 10229 6273 10232 6307
rect 10183 6267 10232 6273
rect 10060 6236 10088 6267
rect 10226 6264 10232 6267
rect 10284 6264 10290 6316
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10888 6304 10916 6344
rect 11333 6341 11345 6344
rect 11379 6341 11391 6375
rect 11333 6335 11391 6341
rect 12250 6332 12256 6384
rect 12308 6332 12314 6384
rect 12710 6332 12716 6384
rect 12768 6332 12774 6384
rect 14182 6332 14188 6384
rect 14240 6332 14246 6384
rect 14734 6332 14740 6384
rect 14792 6372 14798 6384
rect 15197 6375 15255 6381
rect 15197 6372 15209 6375
rect 14792 6344 15209 6372
rect 14792 6332 14798 6344
rect 15197 6341 15209 6344
rect 15243 6372 15255 6375
rect 16040 6372 16068 6412
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 17589 6443 17647 6449
rect 17589 6409 17601 6443
rect 17635 6440 17647 6443
rect 17862 6440 17868 6452
rect 17635 6412 17868 6440
rect 17635 6409 17647 6412
rect 17589 6403 17647 6409
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19518 6440 19524 6452
rect 19392 6412 19524 6440
rect 19392 6400 19398 6412
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 19702 6400 19708 6452
rect 19760 6440 19766 6452
rect 20717 6443 20775 6449
rect 20717 6440 20729 6443
rect 19760 6412 20729 6440
rect 19760 6400 19766 6412
rect 20717 6409 20729 6412
rect 20763 6409 20775 6443
rect 20717 6403 20775 6409
rect 22747 6443 22805 6449
rect 22747 6409 22759 6443
rect 22793 6440 22805 6443
rect 22793 6412 23060 6440
rect 22793 6409 22805 6412
rect 22747 6403 22805 6409
rect 19978 6372 19984 6384
rect 15243 6344 16068 6372
rect 15243 6341 15255 6344
rect 15197 6335 15255 6341
rect 10459 6276 10916 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11020 6276 11529 6304
rect 11020 6264 11026 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 12434 6264 12440 6316
rect 12492 6264 12498 6316
rect 12894 6264 12900 6316
rect 12952 6264 12958 6316
rect 13262 6264 13268 6316
rect 13320 6264 13326 6316
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6304 14979 6307
rect 15010 6304 15016 6316
rect 14967 6276 15016 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6273 15163 6307
rect 15105 6267 15163 6273
rect 10318 6236 10324 6248
rect 10060 6208 10324 6236
rect 10318 6196 10324 6208
rect 10376 6236 10382 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 10376 6208 10517 6236
rect 10376 6196 10382 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 11054 6236 11060 6248
rect 10836 6208 11060 6236
rect 10836 6196 10842 6208
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11606 6196 11612 6248
rect 11664 6236 11670 6248
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 11664 6208 12633 6236
rect 11664 6196 11670 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 10042 6168 10048 6180
rect 9876 6140 10048 6168
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 15120 6168 15148 6267
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 15930 6304 15936 6316
rect 15528 6276 15936 6304
rect 15528 6264 15534 6276
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16040 6313 16068 6344
rect 19444 6344 19984 6372
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16853 6307 16911 6313
rect 16356 6276 16401 6304
rect 16356 6264 16362 6276
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 16942 6304 16948 6316
rect 16899 6276 16948 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6304 17187 6307
rect 17218 6304 17224 6316
rect 17175 6276 17224 6304
rect 17175 6273 17187 6276
rect 17129 6267 17187 6273
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 18138 6304 18144 6316
rect 17543 6276 18144 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 19242 6264 19248 6316
rect 19300 6264 19306 6316
rect 19444 6313 19472 6344
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 20349 6375 20407 6381
rect 20349 6341 20361 6375
rect 20395 6372 20407 6375
rect 20809 6375 20867 6381
rect 20809 6372 20821 6375
rect 20395 6344 20821 6372
rect 20395 6341 20407 6344
rect 20349 6335 20407 6341
rect 20809 6341 20821 6344
rect 20855 6341 20867 6375
rect 20809 6335 20867 6341
rect 21836 6344 22508 6372
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 19518 6264 19524 6316
rect 19576 6264 19582 6316
rect 19702 6264 19708 6316
rect 19760 6264 19766 6316
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 15286 6196 15292 6248
rect 15344 6196 15350 6248
rect 15838 6196 15844 6248
rect 15896 6236 15902 6248
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 15896 6208 16129 6236
rect 15896 6196 15902 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 17034 6236 17040 6248
rect 16117 6199 16175 6205
rect 16224 6208 17040 6236
rect 16224 6168 16252 6208
rect 17034 6196 17040 6208
rect 17092 6196 17098 6248
rect 19058 6196 19064 6248
rect 19116 6236 19122 6248
rect 19720 6236 19748 6264
rect 19116 6208 19748 6236
rect 19116 6196 19122 6208
rect 16945 6171 17003 6177
rect 16945 6168 16957 6171
rect 15120 6140 16252 6168
rect 16500 6140 16957 6168
rect 11330 6100 11336 6112
rect 9784 6072 11336 6100
rect 11330 6060 11336 6072
rect 11388 6100 11394 6112
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 11388 6072 12541 6100
rect 11388 6060 11394 6072
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 12529 6063 12587 6069
rect 14366 6060 14372 6112
rect 14424 6100 14430 6112
rect 14691 6103 14749 6109
rect 14691 6100 14703 6103
rect 14424 6072 14703 6100
rect 14424 6060 14430 6072
rect 14691 6069 14703 6072
rect 14737 6069 14749 6103
rect 14691 6063 14749 6069
rect 15102 6060 15108 6112
rect 15160 6100 15166 6112
rect 15672 6109 15700 6140
rect 15197 6103 15255 6109
rect 15197 6100 15209 6103
rect 15160 6072 15209 6100
rect 15160 6060 15166 6072
rect 15197 6069 15209 6072
rect 15243 6069 15255 6103
rect 15197 6063 15255 6069
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6069 15715 6103
rect 15657 6063 15715 6069
rect 15838 6060 15844 6112
rect 15896 6060 15902 6112
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 16500 6100 16528 6140
rect 16945 6137 16957 6140
rect 16991 6168 17003 6171
rect 17954 6168 17960 6180
rect 16991 6140 17960 6168
rect 16991 6137 17003 6140
rect 16945 6131 17003 6137
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 19334 6128 19340 6180
rect 19392 6128 19398 6180
rect 19812 6112 19840 6267
rect 20162 6264 20168 6316
rect 20220 6264 20226 6316
rect 20438 6264 20444 6316
rect 20496 6264 20502 6316
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 20346 6196 20352 6248
rect 20404 6236 20410 6248
rect 20548 6236 20576 6267
rect 20990 6264 20996 6316
rect 21048 6264 21054 6316
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6273 21235 6307
rect 21177 6267 21235 6273
rect 20404 6208 20576 6236
rect 20404 6196 20410 6208
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 21192 6236 21220 6267
rect 21266 6264 21272 6316
rect 21324 6264 21330 6316
rect 21836 6313 21864 6344
rect 21821 6307 21879 6313
rect 21821 6273 21833 6307
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6304 22063 6307
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 22051 6276 22293 6304
rect 22051 6273 22063 6276
rect 22005 6267 22063 6273
rect 22281 6273 22293 6276
rect 22327 6304 22339 6307
rect 22370 6304 22376 6316
rect 22327 6276 22376 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 22370 6264 22376 6276
rect 22428 6264 22434 6316
rect 22480 6313 22508 6344
rect 22465 6307 22523 6313
rect 22465 6273 22477 6307
rect 22511 6304 22523 6307
rect 22554 6304 22560 6316
rect 22511 6276 22560 6304
rect 22511 6273 22523 6276
rect 22465 6267 22523 6273
rect 22554 6264 22560 6276
rect 22612 6264 22618 6316
rect 22646 6264 22652 6316
rect 22704 6264 22710 6316
rect 22738 6264 22744 6316
rect 22796 6304 22802 6316
rect 22833 6307 22891 6313
rect 22833 6304 22845 6307
rect 22796 6276 22845 6304
rect 22796 6264 22802 6276
rect 22833 6273 22845 6276
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 22922 6264 22928 6316
rect 22980 6264 22986 6316
rect 23032 6304 23060 6412
rect 24118 6332 24124 6384
rect 24176 6332 24182 6384
rect 23385 6307 23443 6313
rect 23385 6304 23397 6307
rect 23032 6276 23397 6304
rect 23385 6273 23397 6276
rect 23431 6273 23443 6307
rect 23385 6267 23443 6273
rect 20680 6208 21220 6236
rect 20680 6196 20686 6208
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 23017 6239 23075 6245
rect 23017 6236 23029 6239
rect 21968 6208 23029 6236
rect 21968 6196 21974 6208
rect 23017 6205 23029 6208
rect 23063 6205 23075 6239
rect 23017 6199 23075 6205
rect 15988 6072 16528 6100
rect 15988 6060 15994 6072
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 16669 6103 16727 6109
rect 16669 6100 16681 6103
rect 16632 6072 16681 6100
rect 16632 6060 16638 6072
rect 16669 6069 16681 6072
rect 16715 6069 16727 6103
rect 16669 6063 16727 6069
rect 19702 6060 19708 6112
rect 19760 6060 19766 6112
rect 19794 6060 19800 6112
rect 19852 6060 19858 6112
rect 19978 6060 19984 6112
rect 20036 6060 20042 6112
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 22189 6103 22247 6109
rect 22189 6100 22201 6103
rect 22060 6072 22201 6100
rect 22060 6060 22066 6072
rect 22189 6069 22201 6072
rect 22235 6069 22247 6103
rect 22189 6063 22247 6069
rect 22278 6060 22284 6112
rect 22336 6060 22342 6112
rect 22370 6060 22376 6112
rect 22428 6100 22434 6112
rect 24811 6103 24869 6109
rect 24811 6100 24823 6103
rect 22428 6072 24823 6100
rect 22428 6060 22434 6072
rect 24811 6069 24823 6072
rect 24857 6069 24869 6103
rect 24811 6063 24869 6069
rect 1104 6010 26312 6032
rect 1104 5958 4101 6010
rect 4153 5958 4165 6010
rect 4217 5958 4229 6010
rect 4281 5958 4293 6010
rect 4345 5958 4357 6010
rect 4409 5958 10403 6010
rect 10455 5958 10467 6010
rect 10519 5958 10531 6010
rect 10583 5958 10595 6010
rect 10647 5958 10659 6010
rect 10711 5958 16705 6010
rect 16757 5958 16769 6010
rect 16821 5958 16833 6010
rect 16885 5958 16897 6010
rect 16949 5958 16961 6010
rect 17013 5958 23007 6010
rect 23059 5958 23071 6010
rect 23123 5958 23135 6010
rect 23187 5958 23199 6010
rect 23251 5958 23263 6010
rect 23315 5958 26312 6010
rect 1104 5936 26312 5958
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 6733 5899 6791 5905
rect 6733 5896 6745 5899
rect 3844 5868 6745 5896
rect 3844 5856 3850 5868
rect 6733 5865 6745 5868
rect 6779 5896 6791 5899
rect 8110 5896 8116 5908
rect 6779 5868 8116 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 9769 5899 9827 5905
rect 8220 5868 9720 5896
rect 6178 5788 6184 5840
rect 6236 5828 6242 5840
rect 7190 5828 7196 5840
rect 6236 5800 7196 5828
rect 6236 5788 6242 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 7469 5831 7527 5837
rect 7469 5797 7481 5831
rect 7515 5797 7527 5831
rect 7469 5791 7527 5797
rect 7098 5720 7104 5772
rect 7156 5720 7162 5772
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6822 5692 6828 5704
rect 6052 5664 6828 5692
rect 6052 5652 6058 5664
rect 6822 5652 6828 5664
rect 6880 5692 6886 5704
rect 7484 5692 7512 5791
rect 7558 5788 7564 5840
rect 7616 5788 7622 5840
rect 7650 5720 7656 5772
rect 7708 5720 7714 5772
rect 8220 5760 8248 5868
rect 8570 5788 8576 5840
rect 8628 5788 8634 5840
rect 9582 5828 9588 5840
rect 8680 5800 9588 5828
rect 7760 5732 8248 5760
rect 7760 5692 7788 5732
rect 8294 5720 8300 5772
rect 8352 5720 8358 5772
rect 6880 5664 7788 5692
rect 6880 5652 6886 5664
rect 7834 5652 7840 5704
rect 7892 5652 7898 5704
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 8680 5624 8708 5800
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 8757 5763 8815 5769
rect 8757 5729 8769 5763
rect 8803 5729 8815 5763
rect 8757 5723 8815 5729
rect 8772 5692 8800 5723
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9692 5760 9720 5868
rect 9769 5865 9781 5899
rect 9815 5896 9827 5899
rect 9950 5896 9956 5908
rect 9815 5868 9956 5896
rect 9815 5865 9827 5868
rect 9769 5859 9827 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 10042 5856 10048 5908
rect 10100 5856 10106 5908
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 11112 5868 12817 5896
rect 11112 5856 11118 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 14182 5856 14188 5908
rect 14240 5856 14246 5908
rect 14734 5856 14740 5908
rect 14792 5856 14798 5908
rect 15013 5899 15071 5905
rect 15013 5865 15025 5899
rect 15059 5896 15071 5899
rect 15562 5896 15568 5908
rect 15059 5868 15568 5896
rect 15059 5865 15071 5868
rect 15013 5859 15071 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 17126 5856 17132 5908
rect 17184 5896 17190 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17184 5868 17693 5896
rect 17184 5856 17190 5868
rect 17681 5865 17693 5868
rect 17727 5896 17739 5899
rect 18598 5896 18604 5908
rect 17727 5868 18604 5896
rect 17727 5865 17739 5868
rect 17681 5859 17739 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 20441 5899 20499 5905
rect 20441 5865 20453 5899
rect 20487 5896 20499 5899
rect 20622 5896 20628 5908
rect 20487 5868 20628 5896
rect 20487 5865 20499 5868
rect 20441 5859 20499 5865
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 20901 5899 20959 5905
rect 20901 5865 20913 5899
rect 20947 5896 20959 5899
rect 21634 5896 21640 5908
rect 20947 5868 21640 5896
rect 20947 5865 20959 5868
rect 20901 5859 20959 5865
rect 10778 5788 10784 5840
rect 10836 5788 10842 5840
rect 11330 5788 11336 5840
rect 11388 5788 11394 5840
rect 14090 5788 14096 5840
rect 14148 5828 14154 5840
rect 14752 5828 14780 5856
rect 17865 5831 17923 5837
rect 17865 5828 17877 5831
rect 14148 5800 14780 5828
rect 15212 5800 17877 5828
rect 14148 5788 14154 5800
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 8904 5732 9260 5760
rect 8904 5720 8910 5732
rect 9232 5701 9260 5732
rect 9692 5732 10517 5760
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8772 5664 9137 5692
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9218 5695 9276 5701
rect 9218 5661 9230 5695
rect 9264 5661 9276 5695
rect 9218 5655 9276 5661
rect 9590 5695 9648 5701
rect 9590 5661 9602 5695
rect 9636 5694 9648 5695
rect 9692 5694 9720 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 12860 5732 14136 5760
rect 12860 5720 12866 5732
rect 9636 5666 9720 5694
rect 9636 5661 9648 5666
rect 9590 5655 9648 5661
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10226 5692 10232 5704
rect 9824 5664 10232 5692
rect 9824 5652 9830 5664
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10318 5652 10324 5704
rect 10376 5652 10382 5704
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10778 5692 10784 5704
rect 10643 5664 10784 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 6144 5596 8708 5624
rect 6144 5584 6150 5596
rect 8754 5584 8760 5636
rect 8812 5624 8818 5636
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 8812 5596 9413 5624
rect 8812 5584 8818 5596
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9401 5587 9459 5593
rect 9493 5627 9551 5633
rect 9493 5593 9505 5627
rect 9539 5624 9551 5627
rect 10612 5624 10640 5655
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5692 11483 5695
rect 12894 5692 12900 5704
rect 11471 5664 12900 5692
rect 11471 5661 11483 5664
rect 11425 5655 11483 5661
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 14108 5701 14136 5732
rect 15212 5701 15240 5800
rect 17865 5797 17877 5800
rect 17911 5797 17923 5831
rect 17865 5791 17923 5797
rect 19518 5788 19524 5840
rect 19576 5828 19582 5840
rect 20916 5828 20944 5859
rect 21634 5856 21640 5868
rect 21692 5856 21698 5908
rect 22281 5899 22339 5905
rect 22281 5865 22293 5899
rect 22327 5896 22339 5899
rect 22922 5896 22928 5908
rect 22327 5868 22928 5896
rect 22327 5865 22339 5868
rect 22281 5859 22339 5865
rect 22922 5856 22928 5868
rect 22980 5856 22986 5908
rect 19576 5800 20944 5828
rect 25041 5831 25099 5837
rect 19576 5788 19582 5800
rect 25041 5797 25053 5831
rect 25087 5797 25099 5831
rect 25041 5791 25099 5797
rect 15838 5760 15844 5772
rect 15488 5732 15844 5760
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5692 15255 5695
rect 15286 5692 15292 5704
rect 15243 5664 15292 5692
rect 15243 5661 15255 5664
rect 15197 5655 15255 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 15378 5652 15384 5704
rect 15436 5652 15442 5704
rect 15488 5701 15516 5732
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 17405 5763 17463 5769
rect 17405 5729 17417 5763
rect 17451 5760 17463 5763
rect 17770 5760 17776 5772
rect 17451 5732 17776 5760
rect 17451 5729 17463 5732
rect 17405 5723 17463 5729
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 21910 5720 21916 5772
rect 21968 5760 21974 5772
rect 22373 5763 22431 5769
rect 22373 5760 22385 5763
rect 21968 5732 22385 5760
rect 21968 5720 21974 5732
rect 22373 5729 22385 5732
rect 22419 5729 22431 5763
rect 22373 5723 22431 5729
rect 22554 5720 22560 5772
rect 22612 5760 22618 5772
rect 25056 5760 25084 5791
rect 22612 5732 25084 5760
rect 22612 5720 22618 5732
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 15654 5652 15660 5704
rect 15712 5652 15718 5704
rect 17954 5652 17960 5704
rect 18012 5652 18018 5704
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 20312 5664 20361 5692
rect 20312 5652 20318 5664
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 20349 5655 20407 5661
rect 22097 5695 22155 5701
rect 22097 5661 22109 5695
rect 22143 5692 22155 5695
rect 22278 5692 22284 5704
rect 22143 5664 22284 5692
rect 22143 5661 22155 5664
rect 22097 5655 22155 5661
rect 9539 5596 10640 5624
rect 10965 5627 11023 5633
rect 9539 5593 9551 5596
rect 9493 5587 9551 5593
rect 10965 5593 10977 5627
rect 11011 5624 11023 5627
rect 11692 5627 11750 5633
rect 11011 5596 11652 5624
rect 11011 5593 11023 5596
rect 10965 5587 11023 5593
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 8021 5559 8079 5565
rect 8021 5556 8033 5559
rect 7708 5528 8033 5556
rect 7708 5516 7714 5528
rect 8021 5525 8033 5528
rect 8067 5525 8079 5559
rect 8021 5519 8079 5525
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 11054 5556 11060 5568
rect 8352 5528 11060 5556
rect 8352 5516 8358 5528
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 11514 5556 11520 5568
rect 11195 5528 11520 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11624 5556 11652 5596
rect 11692 5593 11704 5627
rect 11738 5624 11750 5627
rect 13170 5624 13176 5636
rect 11738 5596 13176 5624
rect 11738 5593 11750 5596
rect 11692 5587 11750 5593
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 14553 5627 14611 5633
rect 14553 5593 14565 5627
rect 14599 5624 14611 5627
rect 15396 5624 15424 5652
rect 14599 5596 15424 5624
rect 14599 5593 14611 5596
rect 14553 5587 14611 5593
rect 17218 5584 17224 5636
rect 17276 5624 17282 5636
rect 17497 5627 17555 5633
rect 17497 5624 17509 5627
rect 17276 5596 17509 5624
rect 17276 5584 17282 5596
rect 17497 5593 17509 5596
rect 17543 5593 17555 5627
rect 17497 5587 17555 5593
rect 11974 5556 11980 5568
rect 11624 5528 11980 5556
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 14734 5516 14740 5568
rect 14792 5565 14798 5568
rect 14792 5559 14811 5565
rect 14799 5525 14811 5559
rect 14792 5519 14811 5525
rect 14792 5516 14798 5519
rect 14918 5516 14924 5568
rect 14976 5516 14982 5568
rect 15381 5559 15439 5565
rect 15381 5525 15393 5559
rect 15427 5556 15439 5559
rect 16390 5556 16396 5568
rect 15427 5528 16396 5556
rect 15427 5525 15439 5528
rect 15381 5519 15439 5525
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 17697 5559 17755 5565
rect 17697 5556 17709 5559
rect 16724 5528 17709 5556
rect 16724 5516 16730 5528
rect 17697 5525 17709 5528
rect 17743 5525 17755 5559
rect 17697 5519 17755 5525
rect 18046 5516 18052 5568
rect 18104 5516 18110 5568
rect 20364 5556 20392 5655
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 22738 5652 22744 5704
rect 22796 5652 22802 5704
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 20717 5627 20775 5633
rect 20717 5593 20729 5627
rect 20763 5624 20775 5627
rect 20806 5624 20812 5636
rect 20763 5596 20812 5624
rect 20763 5593 20775 5596
rect 20717 5587 20775 5593
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 20933 5627 20991 5633
rect 20933 5593 20945 5627
rect 20979 5624 20991 5627
rect 21726 5624 21732 5636
rect 20979 5596 21732 5624
rect 20979 5593 20991 5596
rect 20933 5587 20991 5593
rect 21726 5584 21732 5596
rect 21784 5624 21790 5636
rect 21913 5627 21971 5633
rect 21913 5624 21925 5627
rect 21784 5596 21925 5624
rect 21784 5584 21790 5596
rect 21913 5593 21925 5596
rect 21959 5624 21971 5627
rect 22002 5624 22008 5636
rect 21959 5596 22008 5624
rect 21959 5593 21971 5596
rect 21913 5587 21971 5593
rect 22002 5584 22008 5596
rect 22060 5584 22066 5636
rect 23566 5584 23572 5636
rect 23624 5584 23630 5636
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 20364 5528 21097 5556
rect 21085 5525 21097 5528
rect 21131 5525 21143 5559
rect 21085 5519 21143 5525
rect 22370 5516 22376 5568
rect 22428 5556 22434 5568
rect 24167 5559 24225 5565
rect 24167 5556 24179 5559
rect 22428 5528 24179 5556
rect 22428 5516 22434 5528
rect 24167 5525 24179 5528
rect 24213 5556 24225 5559
rect 24872 5556 24900 5655
rect 24213 5528 24900 5556
rect 24213 5525 24225 5528
rect 24167 5519 24225 5525
rect 1104 5466 26312 5488
rect 1104 5414 4761 5466
rect 4813 5414 4825 5466
rect 4877 5414 4889 5466
rect 4941 5414 4953 5466
rect 5005 5414 5017 5466
rect 5069 5414 11063 5466
rect 11115 5414 11127 5466
rect 11179 5414 11191 5466
rect 11243 5414 11255 5466
rect 11307 5414 11319 5466
rect 11371 5414 17365 5466
rect 17417 5414 17429 5466
rect 17481 5414 17493 5466
rect 17545 5414 17557 5466
rect 17609 5414 17621 5466
rect 17673 5414 23667 5466
rect 23719 5414 23731 5466
rect 23783 5414 23795 5466
rect 23847 5414 23859 5466
rect 23911 5414 23923 5466
rect 23975 5414 26312 5466
rect 1104 5392 26312 5414
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5776 5324 6377 5352
rect 5776 5312 5782 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 7190 5312 7196 5364
rect 7248 5361 7254 5364
rect 7248 5355 7267 5361
rect 7255 5352 7267 5355
rect 7653 5355 7711 5361
rect 7255 5324 7512 5352
rect 7255 5321 7267 5324
rect 7248 5315 7267 5321
rect 7248 5312 7254 5315
rect 6730 5284 6736 5296
rect 6564 5256 6736 5284
rect 6564 5225 6592 5256
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 7009 5287 7067 5293
rect 7009 5253 7021 5287
rect 7055 5253 7067 5287
rect 7009 5247 7067 5253
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 6914 5176 6920 5228
rect 6972 5176 6978 5228
rect 6822 5108 6828 5160
rect 6880 5108 6886 5160
rect 7024 5148 7052 5247
rect 7484 5225 7512 5324
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 7834 5352 7840 5364
rect 7699 5324 7840 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 11606 5352 11612 5364
rect 10275 5324 11612 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15252 5324 15577 5352
rect 15252 5312 15258 5324
rect 15565 5321 15577 5324
rect 15611 5321 15623 5355
rect 15565 5315 15623 5321
rect 16390 5312 16396 5364
rect 16448 5312 16454 5364
rect 16482 5312 16488 5364
rect 16540 5352 16546 5364
rect 16761 5355 16819 5361
rect 16761 5352 16773 5355
rect 16540 5324 16773 5352
rect 16540 5312 16546 5324
rect 16761 5321 16773 5324
rect 16807 5321 16819 5355
rect 17218 5352 17224 5364
rect 16761 5315 16819 5321
rect 16960 5324 17224 5352
rect 15102 5284 15108 5296
rect 14292 5256 15108 5284
rect 14292 5228 14320 5256
rect 15102 5244 15108 5256
rect 15160 5244 15166 5296
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7616 5188 7665 5216
rect 7616 5176 7622 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 7760 5148 7788 5179
rect 7834 5176 7840 5228
rect 7892 5176 7898 5228
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10376 5188 10425 5216
rect 10376 5176 10382 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 14274 5176 14280 5228
rect 14332 5176 14338 5228
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 14976 5188 15761 5216
rect 14976 5176 14982 5188
rect 15749 5185 15761 5188
rect 15795 5216 15807 5219
rect 16301 5219 16359 5225
rect 16301 5216 16313 5219
rect 15795 5188 16313 5216
rect 15795 5185 15807 5188
rect 15749 5179 15807 5185
rect 16301 5185 16313 5188
rect 16347 5185 16359 5219
rect 16408 5216 16436 5312
rect 16960 5225 16988 5324
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 20254 5352 20260 5364
rect 20312 5361 20318 5364
rect 20312 5355 20336 5361
rect 19552 5324 20260 5352
rect 19552 5296 19580 5324
rect 20254 5312 20260 5324
rect 20324 5321 20336 5355
rect 20312 5315 20336 5321
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5352 20499 5355
rect 20990 5352 20996 5364
rect 20487 5324 20996 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 20312 5312 20318 5315
rect 20990 5312 20996 5324
rect 21048 5352 21054 5364
rect 22373 5355 22431 5361
rect 21048 5324 22140 5352
rect 21048 5312 21054 5324
rect 17126 5244 17132 5296
rect 17184 5244 17190 5296
rect 18046 5284 18052 5296
rect 17344 5256 18052 5284
rect 16945 5219 17003 5225
rect 16408 5188 16712 5216
rect 16301 5179 16359 5185
rect 9490 5148 9496 5160
rect 7024 5120 9496 5148
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 10778 5148 10784 5160
rect 10735 5120 10784 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 10778 5108 10784 5120
rect 10836 5148 10842 5160
rect 11054 5148 11060 5160
rect 10836 5120 11060 5148
rect 10836 5108 10842 5120
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 14093 5151 14151 5157
rect 14093 5117 14105 5151
rect 14139 5148 14151 5151
rect 14366 5148 14372 5160
rect 14139 5120 14372 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 7377 5083 7435 5089
rect 7377 5049 7389 5083
rect 7423 5080 7435 5083
rect 7926 5080 7932 5092
rect 7423 5052 7932 5080
rect 7423 5049 7435 5052
rect 7377 5043 7435 5049
rect 7926 5040 7932 5052
rect 7984 5040 7990 5092
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 7064 4984 7205 5012
rect 7064 4972 7070 4984
rect 7193 4981 7205 4984
rect 7239 5012 7251 5015
rect 7558 5012 7564 5024
rect 7239 4984 7564 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10962 5012 10968 5024
rect 10643 4984 10968 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11146 4972 11152 5024
rect 11204 5012 11210 5024
rect 11606 5012 11612 5024
rect 11204 4984 11612 5012
rect 11204 4972 11210 4984
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 14240 4984 14473 5012
rect 14240 4972 14246 4984
rect 14461 4981 14473 4984
rect 14507 5012 14519 5015
rect 14734 5012 14740 5024
rect 14507 4984 14740 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 14734 4972 14740 4984
rect 14792 5012 14798 5024
rect 14918 5012 14924 5024
rect 14792 4984 14924 5012
rect 14792 4972 14798 4984
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15764 5012 15792 5179
rect 15838 5108 15844 5160
rect 15896 5108 15902 5160
rect 15930 5108 15936 5160
rect 15988 5108 15994 5160
rect 16025 5151 16083 5157
rect 16025 5117 16037 5151
rect 16071 5148 16083 5151
rect 16574 5148 16580 5160
rect 16071 5120 16580 5148
rect 16071 5117 16083 5120
rect 16025 5111 16083 5117
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 16684 5148 16712 5188
rect 16945 5185 16957 5219
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17144 5216 17172 5244
rect 17083 5188 17172 5216
rect 17221 5219 17279 5225
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17221 5185 17233 5219
rect 17267 5216 17279 5219
rect 17344 5216 17372 5256
rect 18046 5244 18052 5256
rect 18104 5244 18110 5296
rect 19337 5287 19395 5293
rect 19337 5253 19349 5287
rect 19383 5284 19395 5287
rect 19426 5284 19432 5296
rect 19383 5256 19432 5284
rect 19383 5253 19395 5256
rect 19337 5247 19395 5253
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 19518 5244 19524 5296
rect 19576 5293 19582 5296
rect 19576 5287 19595 5293
rect 19583 5253 19595 5287
rect 19576 5247 19595 5253
rect 19576 5244 19582 5247
rect 19978 5244 19984 5296
rect 20036 5284 20042 5296
rect 20073 5287 20131 5293
rect 20073 5284 20085 5287
rect 20036 5256 20085 5284
rect 20036 5244 20042 5256
rect 20073 5253 20085 5256
rect 20119 5253 20131 5287
rect 20073 5247 20131 5253
rect 17267 5188 17372 5216
rect 17267 5185 17279 5188
rect 17221 5179 17279 5185
rect 17402 5176 17408 5228
rect 17460 5176 17466 5228
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 22112 5216 22140 5324
rect 22373 5321 22385 5355
rect 22419 5352 22431 5355
rect 22738 5352 22744 5364
rect 22419 5324 22744 5352
rect 22419 5321 22431 5324
rect 22373 5315 22431 5321
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 22480 5256 22876 5284
rect 22480 5225 22508 5256
rect 22848 5228 22876 5256
rect 22281 5219 22339 5225
rect 22281 5216 22293 5219
rect 22060 5188 22293 5216
rect 22060 5176 22066 5188
rect 22281 5185 22293 5188
rect 22327 5185 22339 5219
rect 22281 5179 22339 5185
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 17681 5151 17739 5157
rect 17681 5148 17693 5151
rect 16684 5120 17693 5148
rect 17681 5117 17693 5120
rect 17727 5117 17739 5151
rect 17681 5111 17739 5117
rect 20438 5108 20444 5160
rect 20496 5148 20502 5160
rect 22480 5148 22508 5179
rect 22554 5176 22560 5228
rect 22612 5216 22618 5228
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 22612 5188 22661 5216
rect 22612 5176 22618 5188
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 22830 5176 22836 5228
rect 22888 5176 22894 5228
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 20496 5120 22508 5148
rect 20496 5108 20502 5120
rect 16206 5040 16212 5092
rect 16264 5080 16270 5092
rect 17034 5080 17040 5092
rect 16264 5052 17040 5080
rect 16264 5040 16270 5052
rect 17034 5040 17040 5052
rect 17092 5080 17098 5092
rect 17129 5083 17187 5089
rect 17129 5080 17141 5083
rect 17092 5052 17141 5080
rect 17092 5040 17098 5052
rect 17129 5049 17141 5052
rect 17175 5049 17187 5083
rect 17129 5043 17187 5049
rect 19628 5052 20300 5080
rect 19628 5024 19656 5052
rect 16574 5012 16580 5024
rect 15764 4984 16580 5012
rect 16574 4972 16580 4984
rect 16632 5012 16638 5024
rect 16666 5012 16672 5024
rect 16632 4984 16672 5012
rect 16632 4972 16638 4984
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17276 4984 17509 5012
rect 17276 4972 17282 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 17954 4972 17960 5024
rect 18012 4972 18018 5024
rect 19521 5015 19579 5021
rect 19521 4981 19533 5015
rect 19567 5012 19579 5015
rect 19610 5012 19616 5024
rect 19567 4984 19616 5012
rect 19567 4981 19579 4984
rect 19521 4975 19579 4981
rect 19610 4972 19616 4984
rect 19668 4972 19674 5024
rect 19705 5015 19763 5021
rect 19705 4981 19717 5015
rect 19751 5012 19763 5015
rect 20070 5012 20076 5024
rect 19751 4984 20076 5012
rect 19751 4981 19763 4984
rect 19705 4975 19763 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 20272 5021 20300 5052
rect 22646 5040 22652 5092
rect 22704 5040 22710 5092
rect 20257 5015 20315 5021
rect 20257 4981 20269 5015
rect 20303 5012 20315 5015
rect 20806 5012 20812 5024
rect 20303 4984 20812 5012
rect 20303 4981 20315 4984
rect 20257 4975 20315 4981
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 1104 4922 26312 4944
rect 1104 4870 4101 4922
rect 4153 4870 4165 4922
rect 4217 4870 4229 4922
rect 4281 4870 4293 4922
rect 4345 4870 4357 4922
rect 4409 4870 10403 4922
rect 10455 4870 10467 4922
rect 10519 4870 10531 4922
rect 10583 4870 10595 4922
rect 10647 4870 10659 4922
rect 10711 4870 16705 4922
rect 16757 4870 16769 4922
rect 16821 4870 16833 4922
rect 16885 4870 16897 4922
rect 16949 4870 16961 4922
rect 17013 4870 23007 4922
rect 23059 4870 23071 4922
rect 23123 4870 23135 4922
rect 23187 4870 23199 4922
rect 23251 4870 23263 4922
rect 23315 4870 26312 4922
rect 1104 4848 26312 4870
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 7834 4808 7840 4820
rect 6236 4780 7840 4808
rect 6236 4768 6242 4780
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 10962 4768 10968 4820
rect 11020 4768 11026 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 11112 4780 12081 4808
rect 11112 4768 11118 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 25961 4811 26019 4817
rect 25961 4808 25973 4811
rect 12069 4771 12127 4777
rect 12406 4780 25973 4808
rect 6365 4743 6423 4749
rect 6365 4709 6377 4743
rect 6411 4709 6423 4743
rect 11514 4740 11520 4752
rect 6365 4703 6423 4709
rect 10980 4712 11520 4740
rect 6380 4672 6408 4703
rect 5184 4644 6408 4672
rect 5184 4613 5212 4644
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5592 4576 5641 4604
rect 5592 4564 5598 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 5905 4607 5963 4613
rect 5905 4604 5917 4607
rect 5776 4576 5917 4604
rect 5776 4564 5782 4576
rect 5905 4573 5917 4576
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6144 4576 6469 4604
rect 6144 4564 6150 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 7650 4564 7656 4616
rect 7708 4564 7714 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 7926 4604 7932 4616
rect 7883 4576 7932 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8478 4564 8484 4616
rect 8536 4564 8542 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4604 10931 4607
rect 10980 4604 11008 4712
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 11698 4700 11704 4752
rect 11756 4740 11762 4752
rect 12406 4740 12434 4780
rect 25961 4777 25973 4780
rect 26007 4777 26019 4811
rect 25961 4771 26019 4777
rect 11756 4712 12434 4740
rect 13541 4743 13599 4749
rect 11756 4700 11762 4712
rect 13541 4709 13553 4743
rect 13587 4740 13599 4743
rect 14550 4740 14556 4752
rect 13587 4712 14556 4740
rect 13587 4709 13599 4712
rect 13541 4703 13599 4709
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 18969 4743 19027 4749
rect 18969 4709 18981 4743
rect 19015 4740 19027 4743
rect 19426 4740 19432 4752
rect 19015 4712 19432 4740
rect 19015 4709 19027 4712
rect 18969 4703 19027 4709
rect 19426 4700 19432 4712
rect 19484 4700 19490 4752
rect 20162 4740 20168 4752
rect 19536 4712 20168 4740
rect 11882 4672 11888 4684
rect 11164 4644 11888 4672
rect 10919 4576 11008 4604
rect 10919 4573 10931 4576
rect 10873 4567 10931 4573
rect 11054 4564 11060 4616
rect 11112 4564 11118 4616
rect 11164 4613 11192 4644
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 14921 4675 14979 4681
rect 14921 4672 14933 4675
rect 13832 4644 14933 4672
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 12618 4604 12624 4616
rect 12023 4576 12624 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 5445 4539 5503 4545
rect 5445 4505 5457 4539
rect 5491 4536 5503 4539
rect 5997 4539 6055 4545
rect 5491 4508 5948 4536
rect 5491 4505 5503 4508
rect 5445 4499 5503 4505
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4672 4440 4997 4468
rect 4672 4428 4678 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 4985 4431 5043 4437
rect 5810 4428 5816 4480
rect 5868 4428 5874 4480
rect 5920 4468 5948 4508
rect 5997 4505 6009 4539
rect 6043 4536 6055 4539
rect 6043 4508 7696 4536
rect 6043 4505 6055 4508
rect 5997 4499 6055 4505
rect 7668 4480 7696 4508
rect 10042 4496 10048 4548
rect 10100 4536 10106 4548
rect 11241 4539 11299 4545
rect 11241 4536 11253 4539
rect 10100 4508 11253 4536
rect 10100 4496 10106 4508
rect 11241 4505 11253 4508
rect 11287 4505 11299 4539
rect 11241 4499 11299 4505
rect 6197 4471 6255 4477
rect 6197 4468 6209 4471
rect 5920 4440 6209 4468
rect 6197 4437 6209 4440
rect 6243 4437 6255 4471
rect 6197 4431 6255 4437
rect 6546 4428 6552 4480
rect 6604 4428 6610 4480
rect 7650 4428 7656 4480
rect 7708 4428 7714 4480
rect 7742 4428 7748 4480
rect 7800 4428 7806 4480
rect 8297 4471 8355 4477
rect 8297 4437 8309 4471
rect 8343 4468 8355 4471
rect 8386 4468 8392 4480
rect 8343 4440 8392 4468
rect 8343 4437 8355 4440
rect 8297 4431 8355 4437
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 11348 4468 11376 4567
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 13832 4613 13860 4644
rect 14921 4641 14933 4644
rect 14967 4672 14979 4675
rect 15010 4672 15016 4684
rect 14967 4644 15016 4672
rect 14967 4641 14979 4644
rect 14921 4635 14979 4641
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 19536 4681 19564 4712
rect 20162 4700 20168 4712
rect 20220 4740 20226 4752
rect 20220 4712 21404 4740
rect 20220 4700 20226 4712
rect 19521 4675 19579 4681
rect 19521 4641 19533 4675
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 19610 4632 19616 4684
rect 19668 4672 19674 4684
rect 19668 4644 20116 4672
rect 19668 4632 19674 4644
rect 13817 4607 13875 4613
rect 13817 4573 13829 4607
rect 13863 4573 13875 4607
rect 13817 4567 13875 4573
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14458 4613 14464 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13964 4576 14289 4604
rect 13964 4564 13970 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14455 4567 14464 4613
rect 14516 4604 14522 4616
rect 15197 4607 15255 4613
rect 14516 4576 14555 4604
rect 14458 4564 14464 4567
rect 14516 4564 14522 4576
rect 15197 4573 15209 4607
rect 15243 4604 15255 4607
rect 15286 4604 15292 4616
rect 15243 4576 15292 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 16574 4564 16580 4616
rect 16632 4564 16638 4616
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4604 16819 4607
rect 17402 4604 17408 4616
rect 16807 4576 17408 4604
rect 16807 4573 16819 4576
rect 16761 4567 16819 4573
rect 13541 4539 13599 4545
rect 13541 4505 13553 4539
rect 13587 4536 13599 4539
rect 13630 4536 13636 4548
rect 13587 4508 13636 4536
rect 13587 4505 13599 4508
rect 13541 4499 13599 4505
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 13998 4496 14004 4548
rect 14056 4536 14062 4548
rect 14369 4539 14427 4545
rect 14369 4536 14381 4539
rect 14056 4508 14381 4536
rect 14056 4496 14062 4508
rect 14369 4505 14381 4508
rect 14415 4505 14427 4539
rect 14369 4499 14427 4505
rect 14553 4539 14611 4545
rect 14553 4505 14565 4539
rect 14599 4505 14611 4539
rect 14553 4499 14611 4505
rect 11020 4440 11376 4468
rect 14568 4468 14596 4499
rect 14734 4496 14740 4548
rect 14792 4496 14798 4548
rect 14826 4496 14832 4548
rect 14884 4536 14890 4548
rect 15013 4539 15071 4545
rect 15013 4536 15025 4539
rect 14884 4508 15025 4536
rect 14884 4496 14890 4508
rect 15013 4505 15025 4508
rect 15059 4505 15071 4539
rect 15013 4499 15071 4505
rect 15930 4496 15936 4548
rect 15988 4536 15994 4548
rect 16776 4536 16804 4567
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 15988 4508 16804 4536
rect 18892 4536 18920 4567
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 20088 4613 20116 4644
rect 20254 4632 20260 4684
rect 20312 4632 20318 4684
rect 20438 4632 20444 4684
rect 20496 4672 20502 4684
rect 20533 4675 20591 4681
rect 20533 4672 20545 4675
rect 20496 4644 20545 4672
rect 20496 4632 20502 4644
rect 20533 4641 20545 4644
rect 20579 4641 20591 4675
rect 20533 4635 20591 4641
rect 20806 4632 20812 4684
rect 20864 4632 20870 4684
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 21008 4644 21281 4672
rect 21008 4613 21036 4644
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 19889 4607 19947 4613
rect 19889 4604 19901 4607
rect 19751 4576 19901 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 19889 4573 19901 4576
rect 19935 4573 19947 4607
rect 19889 4567 19947 4573
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4573 20131 4607
rect 20073 4567 20131 4573
rect 20349 4607 20407 4613
rect 20349 4573 20361 4607
rect 20395 4604 20407 4607
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20395 4576 20729 4604
rect 20395 4573 20407 4576
rect 20349 4567 20407 4573
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20717 4567 20775 4573
rect 20824 4576 20913 4604
rect 19978 4536 19984 4548
rect 18892 4508 19984 4536
rect 15988 4496 15994 4508
rect 19978 4496 19984 4508
rect 20036 4536 20042 4548
rect 20364 4536 20392 4567
rect 20036 4508 20392 4536
rect 20036 4496 20042 4508
rect 14918 4468 14924 4480
rect 14568 4440 14924 4468
rect 11020 4428 11026 4440
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15378 4428 15384 4480
rect 15436 4428 15442 4480
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 16945 4471 17003 4477
rect 16945 4468 16957 4471
rect 16908 4440 16957 4468
rect 16908 4428 16914 4440
rect 16945 4437 16957 4440
rect 16991 4437 17003 4471
rect 16945 4431 17003 4437
rect 19242 4428 19248 4480
rect 19300 4428 19306 4480
rect 20254 4428 20260 4480
rect 20312 4468 20318 4480
rect 20824 4468 20852 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 21177 4607 21235 4613
rect 21177 4573 21189 4607
rect 21223 4604 21235 4607
rect 21376 4604 21404 4712
rect 21726 4632 21732 4684
rect 21784 4632 21790 4684
rect 22005 4675 22063 4681
rect 22005 4641 22017 4675
rect 22051 4672 22063 4675
rect 22051 4644 22140 4672
rect 22051 4641 22063 4644
rect 22005 4635 22063 4641
rect 21223 4576 21404 4604
rect 21223 4573 21235 4576
rect 21177 4567 21235 4573
rect 20990 4468 20996 4480
rect 20312 4440 20996 4468
rect 20312 4428 20318 4440
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 21192 4468 21220 4567
rect 21634 4564 21640 4616
rect 21692 4564 21698 4616
rect 22112 4613 22140 4644
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4573 22155 4607
rect 22097 4567 22155 4573
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 22002 4496 22008 4548
rect 22060 4536 22066 4548
rect 22296 4536 22324 4567
rect 25774 4564 25780 4616
rect 25832 4564 25838 4616
rect 22060 4508 22324 4536
rect 22060 4496 22066 4508
rect 22370 4468 22376 4480
rect 21192 4440 22376 4468
rect 22370 4428 22376 4440
rect 22428 4428 22434 4480
rect 22462 4428 22468 4480
rect 22520 4428 22526 4480
rect 1104 4378 26312 4400
rect 1104 4326 4761 4378
rect 4813 4326 4825 4378
rect 4877 4326 4889 4378
rect 4941 4326 4953 4378
rect 5005 4326 5017 4378
rect 5069 4326 11063 4378
rect 11115 4326 11127 4378
rect 11179 4326 11191 4378
rect 11243 4326 11255 4378
rect 11307 4326 11319 4378
rect 11371 4326 17365 4378
rect 17417 4326 17429 4378
rect 17481 4326 17493 4378
rect 17545 4326 17557 4378
rect 17609 4326 17621 4378
rect 17673 4326 23667 4378
rect 23719 4326 23731 4378
rect 23783 4326 23795 4378
rect 23847 4326 23859 4378
rect 23911 4326 23923 4378
rect 23975 4326 26312 4378
rect 1104 4304 26312 4326
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5721 4267 5779 4273
rect 5721 4264 5733 4267
rect 5592 4236 5733 4264
rect 5592 4224 5598 4236
rect 5721 4233 5733 4236
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 5828 4236 7696 4264
rect 4614 4205 4620 4208
rect 4608 4196 4620 4205
rect 4575 4168 4620 4196
rect 4608 4159 4620 4168
rect 4614 4156 4620 4159
rect 4672 4156 4678 4208
rect 5828 4205 5856 4236
rect 7668 4208 7696 4236
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7853 4267 7911 4273
rect 7853 4264 7865 4267
rect 7800 4236 7865 4264
rect 7800 4224 7806 4236
rect 7853 4233 7865 4236
rect 7899 4233 7911 4267
rect 7853 4227 7911 4233
rect 9490 4224 9496 4276
rect 9548 4224 9554 4276
rect 11241 4267 11299 4273
rect 11241 4264 11253 4267
rect 10244 4236 11253 4264
rect 5813 4199 5871 4205
rect 5813 4165 5825 4199
rect 5859 4165 5871 4199
rect 5813 4159 5871 4165
rect 6029 4199 6087 4205
rect 6029 4165 6041 4199
rect 6075 4196 6087 4199
rect 6730 4196 6736 4208
rect 6075 4168 6736 4196
rect 6075 4165 6087 4168
rect 6029 4159 6087 4165
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 7009 4199 7067 4205
rect 7009 4165 7021 4199
rect 7055 4196 7067 4199
rect 7098 4196 7104 4208
rect 7055 4168 7104 4196
rect 7055 4165 7067 4168
rect 7009 4159 7067 4165
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 7209 4199 7267 4205
rect 7209 4196 7221 4199
rect 7208 4165 7221 4196
rect 7255 4165 7267 4199
rect 7208 4159 7267 4165
rect 5626 4128 5632 4140
rect 4356 4100 5632 4128
rect 4356 4069 4384 4100
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 6546 4060 6552 4072
rect 5500 4032 6552 4060
rect 5500 4020 5506 4032
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6656 4060 6684 4091
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7208 4128 7236 4159
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 8202 4196 8208 4208
rect 7708 4168 8208 4196
rect 7708 4156 7714 4168
rect 8202 4156 8208 4168
rect 8260 4196 8266 4208
rect 8260 4168 8524 4196
rect 8260 4156 8266 4168
rect 7926 4128 7932 4140
rect 6963 4100 7932 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 8110 4088 8116 4140
rect 8168 4088 8174 4140
rect 8386 4137 8392 4140
rect 8380 4128 8392 4137
rect 8347 4100 8392 4128
rect 8380 4091 8392 4100
rect 8386 4088 8392 4091
rect 8444 4088 8450 4140
rect 8496 4128 8524 4168
rect 10042 4156 10048 4208
rect 10100 4156 10106 4208
rect 9858 4128 9864 4140
rect 8496 4100 9864 4128
rect 9858 4088 9864 4100
rect 9916 4128 9922 4140
rect 10244 4137 10272 4236
rect 11241 4233 11253 4236
rect 11287 4233 11299 4267
rect 11241 4227 11299 4233
rect 11882 4224 11888 4276
rect 11940 4224 11946 4276
rect 13357 4267 13415 4273
rect 13357 4233 13369 4267
rect 13403 4264 13415 4267
rect 13630 4264 13636 4276
rect 13403 4236 13636 4264
rect 13403 4233 13415 4236
rect 13357 4227 13415 4233
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 13722 4224 13728 4276
rect 13780 4264 13786 4276
rect 14458 4264 14464 4276
rect 13780 4236 14464 4264
rect 13780 4224 13786 4236
rect 14458 4224 14464 4236
rect 14516 4264 14522 4276
rect 16482 4264 16488 4276
rect 14516 4236 16488 4264
rect 14516 4224 14522 4236
rect 16482 4224 16488 4236
rect 16540 4264 16546 4276
rect 17126 4264 17132 4276
rect 16540 4236 17132 4264
rect 16540 4224 16546 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 19978 4224 19984 4276
rect 20036 4264 20042 4276
rect 20073 4267 20131 4273
rect 20073 4264 20085 4267
rect 20036 4236 20085 4264
rect 20036 4224 20042 4236
rect 20073 4233 20085 4236
rect 20119 4233 20131 4267
rect 20073 4227 20131 4233
rect 20806 4224 20812 4276
rect 20864 4224 20870 4276
rect 10778 4196 10784 4208
rect 10612 4168 10784 4196
rect 10612 4137 10640 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 11514 4156 11520 4208
rect 11572 4156 11578 4208
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 11701 4199 11759 4205
rect 11701 4196 11713 4199
rect 11664 4168 11713 4196
rect 11664 4156 11670 4168
rect 11701 4165 11713 4168
rect 11747 4165 11759 4199
rect 11701 4159 11759 4165
rect 14366 4156 14372 4208
rect 14424 4196 14430 4208
rect 16945 4199 17003 4205
rect 14424 4168 14780 4196
rect 14424 4156 14430 4168
rect 10229 4131 10287 4137
rect 10229 4128 10241 4131
rect 9916 4100 10241 4128
rect 9916 4088 9922 4100
rect 10229 4097 10241 4100
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 10962 4128 10968 4140
rect 10597 4091 10655 4097
rect 10704 4100 10968 4128
rect 7098 4060 7104 4072
rect 6656 4032 7104 4060
rect 6932 4004 6960 4032
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 10336 4060 10364 4091
rect 10704 4069 10732 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 11146 4128 11152 4140
rect 11103 4100 11152 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 11333 4131 11391 4137
rect 11333 4097 11345 4131
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 9272 4032 10364 4060
rect 9272 4020 9278 4032
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 5718 3992 5724 4004
rect 5592 3964 5724 3992
rect 5592 3952 5598 3964
rect 5718 3952 5724 3964
rect 5776 3992 5782 4004
rect 6362 3992 6368 4004
rect 5776 3964 6368 3992
rect 5776 3952 5782 3964
rect 6362 3952 6368 3964
rect 6420 3992 6426 4004
rect 6420 3964 6776 3992
rect 6420 3952 6426 3964
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6086 3924 6092 3936
rect 6043 3896 6092 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6178 3884 6184 3936
rect 6236 3884 6242 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6638 3924 6644 3936
rect 6503 3896 6644 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6748 3924 6776 3964
rect 6914 3952 6920 4004
rect 6972 3952 6978 4004
rect 7377 3995 7435 4001
rect 7377 3992 7389 3995
rect 7024 3964 7389 3992
rect 7024 3924 7052 3964
rect 7377 3961 7389 3964
rect 7423 3961 7435 3995
rect 10336 3992 10364 4032
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 11348 4060 11376 4091
rect 11974 4088 11980 4140
rect 12032 4088 12038 4140
rect 12618 4088 12624 4140
rect 12676 4088 12682 4140
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12860 4100 12909 4128
rect 12860 4088 12866 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 10689 4023 10747 4029
rect 10888 4032 11376 4060
rect 10888 3992 10916 4032
rect 10336 3964 10916 3992
rect 10965 3995 11023 4001
rect 7377 3955 7435 3961
rect 10965 3961 10977 3995
rect 11011 3992 11023 3995
rect 11146 3992 11152 4004
rect 11011 3964 11152 3992
rect 11011 3961 11023 3964
rect 10965 3955 11023 3961
rect 11146 3952 11152 3964
rect 11204 3952 11210 4004
rect 13188 3992 13216 4091
rect 14090 4088 14096 4140
rect 14148 4088 14154 4140
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14752 4137 14780 4168
rect 16945 4165 16957 4199
rect 16991 4196 17003 4199
rect 17954 4196 17960 4208
rect 16991 4168 17960 4196
rect 16991 4165 17003 4168
rect 16945 4159 17003 4165
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 19334 4156 19340 4208
rect 19392 4156 19398 4208
rect 20824 4196 20852 4224
rect 20824 4168 21128 4196
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14332 4100 14565 4128
rect 14332 4088 14338 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 15194 4128 15200 4140
rect 15059 4100 15200 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 14182 4020 14188 4072
rect 14240 4020 14246 4072
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4060 14519 4063
rect 14826 4060 14832 4072
rect 14507 4032 14832 4060
rect 14507 4029 14519 4032
rect 14461 4023 14519 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 15028 3992 15056 4091
rect 15194 4088 15200 4100
rect 15252 4128 15258 4140
rect 15838 4128 15844 4140
rect 15252 4100 15844 4128
rect 15252 4088 15258 4100
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15988 4100 16129 4128
rect 15988 4088 15994 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16850 4088 16856 4140
rect 16908 4088 16914 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 16206 4020 16212 4072
rect 16264 4020 16270 4072
rect 17052 4060 17080 4091
rect 17126 4088 17132 4140
rect 17184 4137 17190 4140
rect 17184 4131 17213 4137
rect 17201 4097 17213 4131
rect 17184 4091 17213 4097
rect 17184 4088 17190 4091
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17828 4100 18337 4128
rect 17828 4088 17834 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 20254 4088 20260 4140
rect 20312 4128 20318 4140
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 20312 4100 20453 4128
rect 20312 4088 20318 4100
rect 20441 4097 20453 4100
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 20530 4088 20536 4140
rect 20588 4128 20594 4140
rect 21100 4137 21128 4168
rect 22462 4156 22468 4208
rect 22520 4196 22526 4208
rect 22833 4199 22891 4205
rect 22833 4196 22845 4199
rect 22520 4168 22845 4196
rect 22520 4156 22526 4168
rect 22833 4165 22845 4168
rect 22879 4165 22891 4199
rect 22833 4159 22891 4165
rect 22922 4156 22928 4208
rect 22980 4156 22986 4208
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20588 4100 20821 4128
rect 20588 4088 20594 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 21085 4131 21143 4137
rect 21085 4097 21097 4131
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 21634 4088 21640 4140
rect 21692 4128 21698 4140
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 21692 4100 22201 4128
rect 21692 4088 21698 4100
rect 22189 4097 22201 4100
rect 22235 4128 22247 4131
rect 22370 4128 22376 4140
rect 22235 4100 22376 4128
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22646 4088 22652 4140
rect 22704 4088 22710 4140
rect 23017 4131 23075 4137
rect 23017 4097 23029 4131
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 16408 4032 17080 4060
rect 17313 4063 17371 4069
rect 13188 3964 15056 3992
rect 15565 3995 15623 4001
rect 15565 3961 15577 3995
rect 15611 3992 15623 3995
rect 16408 3992 16436 4032
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4060 18659 4063
rect 19242 4060 19248 4072
rect 18647 4032 19248 4060
rect 18647 4029 18659 4032
rect 18601 4023 18659 4029
rect 15611 3964 16436 3992
rect 16485 3995 16543 4001
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 16485 3961 16497 3995
rect 16531 3992 16543 3995
rect 17328 3992 17356 4023
rect 19242 4020 19248 4032
rect 19300 4020 19306 4072
rect 20070 4020 20076 4072
rect 20128 4060 20134 4072
rect 20349 4063 20407 4069
rect 20349 4060 20361 4063
rect 20128 4032 20361 4060
rect 20128 4020 20134 4032
rect 20349 4029 20361 4032
rect 20395 4029 20407 4063
rect 20349 4023 20407 4029
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 16531 3964 17356 3992
rect 16531 3961 16543 3964
rect 16485 3955 16543 3961
rect 19610 3952 19616 4004
rect 19668 3992 19674 4004
rect 20165 3995 20223 4001
rect 20165 3992 20177 3995
rect 19668 3964 20177 3992
rect 19668 3952 19674 3964
rect 20165 3961 20177 3964
rect 20211 3961 20223 3995
rect 20732 3992 20760 4023
rect 20990 4020 20996 4072
rect 21048 4020 21054 4072
rect 22278 4020 22284 4072
rect 22336 4020 22342 4072
rect 22557 4063 22615 4069
rect 22557 4029 22569 4063
rect 22603 4060 22615 4063
rect 23032 4060 23060 4091
rect 22603 4032 23060 4060
rect 22603 4029 22615 4032
rect 22557 4023 22615 4029
rect 21453 3995 21511 4001
rect 21453 3992 21465 3995
rect 20732 3964 21465 3992
rect 20165 3955 20223 3961
rect 21453 3961 21465 3964
rect 21499 3961 21511 3995
rect 21453 3955 21511 3961
rect 6748 3896 7052 3924
rect 7190 3884 7196 3936
rect 7248 3884 7254 3936
rect 7834 3884 7840 3936
rect 7892 3884 7898 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8478 3924 8484 3936
rect 8067 3896 8484 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 10042 3884 10048 3936
rect 10100 3884 10106 3936
rect 11054 3884 11060 3936
rect 11112 3884 11118 3936
rect 12986 3884 12992 3936
rect 13044 3884 13050 3936
rect 14366 3884 14372 3936
rect 14424 3924 14430 3936
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 14424 3896 14565 3924
rect 14424 3884 14430 3896
rect 14553 3893 14565 3896
rect 14599 3924 14611 3927
rect 14734 3924 14740 3936
rect 14599 3896 14740 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 16669 3927 16727 3933
rect 16669 3893 16681 3927
rect 16715 3924 16727 3927
rect 17034 3924 17040 3936
rect 16715 3896 17040 3924
rect 16715 3893 16727 3896
rect 16669 3887 16727 3893
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 23201 3927 23259 3933
rect 23201 3924 23213 3927
rect 22704 3896 23213 3924
rect 22704 3884 22710 3896
rect 23201 3893 23213 3896
rect 23247 3893 23259 3927
rect 23201 3887 23259 3893
rect 1104 3834 26312 3856
rect 1104 3782 4101 3834
rect 4153 3782 4165 3834
rect 4217 3782 4229 3834
rect 4281 3782 4293 3834
rect 4345 3782 4357 3834
rect 4409 3782 10403 3834
rect 10455 3782 10467 3834
rect 10519 3782 10531 3834
rect 10583 3782 10595 3834
rect 10647 3782 10659 3834
rect 10711 3782 16705 3834
rect 16757 3782 16769 3834
rect 16821 3782 16833 3834
rect 16885 3782 16897 3834
rect 16949 3782 16961 3834
rect 17013 3782 23007 3834
rect 23059 3782 23071 3834
rect 23123 3782 23135 3834
rect 23187 3782 23199 3834
rect 23251 3782 23263 3834
rect 23315 3782 26312 3834
rect 1104 3760 26312 3782
rect 7285 3723 7343 3729
rect 7285 3689 7297 3723
rect 7331 3720 7343 3723
rect 7834 3720 7840 3732
rect 7331 3692 7840 3720
rect 7331 3689 7343 3692
rect 7285 3683 7343 3689
rect 7834 3680 7840 3692
rect 7892 3720 7898 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 7892 3692 8493 3720
rect 7892 3680 7898 3692
rect 8481 3689 8493 3692
rect 8527 3720 8539 3723
rect 9214 3720 9220 3732
rect 8527 3692 9220 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 11793 3723 11851 3729
rect 11793 3689 11805 3723
rect 11839 3720 11851 3723
rect 11974 3720 11980 3732
rect 11839 3692 11980 3720
rect 11839 3689 11851 3692
rect 11793 3683 11851 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 12492 3692 14749 3720
rect 12492 3680 12498 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 14737 3683 14795 3689
rect 17589 3723 17647 3729
rect 17589 3689 17601 3723
rect 17635 3720 17647 3723
rect 18230 3720 18236 3732
rect 17635 3692 18236 3720
rect 17635 3689 17647 3692
rect 17589 3683 17647 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20993 3723 21051 3729
rect 20993 3720 21005 3723
rect 20864 3692 21005 3720
rect 20864 3680 20870 3692
rect 20993 3689 21005 3692
rect 21039 3689 21051 3723
rect 20993 3683 21051 3689
rect 22370 3680 22376 3732
rect 22428 3720 22434 3732
rect 22925 3723 22983 3729
rect 22925 3720 22937 3723
rect 22428 3692 22937 3720
rect 22428 3680 22434 3692
rect 22925 3689 22937 3692
rect 22971 3689 22983 3723
rect 22925 3683 22983 3689
rect 23569 3723 23627 3729
rect 23569 3689 23581 3723
rect 23615 3720 23627 3723
rect 24302 3720 24308 3732
rect 23615 3692 24308 3720
rect 23615 3689 23627 3692
rect 23569 3683 23627 3689
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 7009 3655 7067 3661
rect 7009 3652 7021 3655
rect 6972 3624 7021 3652
rect 6972 3612 6978 3624
rect 7009 3621 7021 3624
rect 7055 3621 7067 3655
rect 8110 3652 8116 3664
rect 7009 3615 7067 3621
rect 7116 3624 8116 3652
rect 5261 3587 5319 3593
rect 5261 3553 5273 3587
rect 5307 3584 5319 3587
rect 5534 3584 5540 3596
rect 5307 3556 5540 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5442 3516 5448 3528
rect 5215 3488 5448 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 7116 3516 7144 3624
rect 8110 3612 8116 3624
rect 8168 3652 8174 3664
rect 8168 3624 8340 3652
rect 8168 3612 8174 3624
rect 7926 3544 7932 3596
rect 7984 3544 7990 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8312 3584 8340 3624
rect 8662 3612 8668 3664
rect 8720 3612 8726 3664
rect 13863 3655 13921 3661
rect 13863 3621 13875 3655
rect 13909 3652 13921 3655
rect 14274 3652 14280 3664
rect 13909 3624 14280 3652
rect 13909 3621 13921 3624
rect 13863 3615 13921 3621
rect 14274 3612 14280 3624
rect 14332 3612 14338 3664
rect 15749 3655 15807 3661
rect 15749 3621 15761 3655
rect 15795 3621 15807 3655
rect 15749 3615 15807 3621
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8312 3556 8953 3584
rect 8205 3547 8263 3553
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 12069 3587 12127 3593
rect 12069 3553 12081 3587
rect 12115 3584 12127 3587
rect 12894 3584 12900 3596
rect 12115 3556 12900 3584
rect 12115 3553 12127 3556
rect 12069 3547 12127 3553
rect 5684 3488 7144 3516
rect 5684 3476 5690 3488
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7248 3488 7849 3516
rect 7248 3476 7254 3488
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 8220 3516 8248 3547
rect 8956 3516 8984 3547
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 14366 3544 14372 3596
rect 14424 3544 14430 3596
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 14691 3556 15608 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 9950 3516 9956 3528
rect 8220 3488 8432 3516
rect 8956 3488 9956 3516
rect 7837 3479 7895 3485
rect 5896 3451 5954 3457
rect 5896 3417 5908 3451
rect 5942 3448 5954 3451
rect 5994 3448 6000 3460
rect 5942 3420 6000 3448
rect 5942 3417 5954 3420
rect 5896 3411 5954 3417
rect 5994 3408 6000 3420
rect 6052 3408 6058 3460
rect 7101 3451 7159 3457
rect 7101 3417 7113 3451
rect 7147 3448 7159 3451
rect 7650 3448 7656 3460
rect 7147 3420 7656 3448
rect 7147 3417 7159 3420
rect 7101 3411 7159 3417
rect 7650 3408 7656 3420
rect 7708 3408 7714 3460
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 4709 3383 4767 3389
rect 4709 3380 4721 3383
rect 4672 3352 4721 3380
rect 4672 3340 4678 3352
rect 4709 3349 4721 3352
rect 4755 3349 4767 3383
rect 4709 3343 4767 3349
rect 5537 3383 5595 3389
rect 5537 3349 5549 3383
rect 5583 3380 5595 3383
rect 7301 3383 7359 3389
rect 7301 3380 7313 3383
rect 5583 3352 7313 3380
rect 5583 3349 5595 3352
rect 5537 3343 5595 3349
rect 7301 3349 7313 3352
rect 7347 3349 7359 3383
rect 7301 3343 7359 3349
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 7852 3380 7880 3479
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 8297 3451 8355 3457
rect 8297 3448 8309 3451
rect 8260 3420 8309 3448
rect 8260 3408 8266 3420
rect 8297 3417 8309 3420
rect 8343 3417 8355 3451
rect 8404 3448 8432 3488
rect 9950 3476 9956 3488
rect 10008 3516 10014 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10008 3488 10425 3516
rect 10008 3476 10014 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10680 3519 10738 3525
rect 10680 3485 10692 3519
rect 10726 3516 10738 3519
rect 11054 3516 11060 3528
rect 10726 3488 11060 3516
rect 10726 3485 10738 3488
rect 10680 3479 10738 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14148 3488 14289 3516
rect 14148 3476 14154 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14608 3488 14749 3516
rect 14608 3476 14614 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 15010 3476 15016 3528
rect 15068 3476 15074 3528
rect 15197 3519 15255 3525
rect 15197 3485 15209 3519
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 8497 3451 8555 3457
rect 8497 3448 8509 3451
rect 8404 3420 8509 3448
rect 8297 3411 8355 3417
rect 8497 3417 8509 3420
rect 8543 3417 8555 3451
rect 8497 3411 8555 3417
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 9186 3451 9244 3457
rect 9186 3448 9198 3451
rect 8812 3420 9198 3448
rect 8812 3408 8818 3420
rect 9186 3417 9198 3420
rect 9232 3417 9244 3451
rect 9186 3411 9244 3417
rect 12986 3408 12992 3460
rect 13044 3408 13050 3460
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 15212 3448 15240 3479
rect 15378 3476 15384 3528
rect 15436 3476 15442 3528
rect 15580 3525 15608 3556
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3485 15623 3519
rect 15764 3516 15792 3615
rect 17770 3612 17776 3664
rect 17828 3612 17834 3664
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3584 15899 3587
rect 17788 3584 17816 3612
rect 19245 3587 19303 3593
rect 19245 3584 19257 3587
rect 15887 3556 19257 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 19245 3553 19257 3556
rect 19291 3584 19303 3587
rect 21177 3587 21235 3593
rect 21177 3584 21189 3587
rect 19291 3556 21189 3584
rect 19291 3553 19303 3556
rect 19245 3547 19303 3553
rect 21177 3553 21189 3556
rect 21223 3553 21235 3587
rect 21177 3547 21235 3553
rect 21545 3587 21603 3593
rect 21545 3553 21557 3587
rect 21591 3584 21603 3587
rect 22646 3584 22652 3596
rect 21591 3556 22652 3584
rect 21591 3553 21603 3556
rect 21545 3547 21603 3553
rect 22646 3544 22652 3556
rect 22704 3544 22710 3596
rect 23584 3584 23612 3683
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 23308 3556 23612 3584
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 15764 3488 16221 3516
rect 15565 3479 15623 3485
rect 16209 3485 16221 3488
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17184 3488 17785 3516
rect 17184 3476 17190 3488
rect 17773 3485 17785 3488
rect 17819 3516 17831 3519
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 17819 3488 18061 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18049 3485 18061 3488
rect 18095 3516 18107 3519
rect 18138 3516 18144 3528
rect 18095 3488 18144 3516
rect 18095 3485 18107 3488
rect 18049 3479 18107 3485
rect 18138 3476 18144 3488
rect 18196 3516 18202 3528
rect 18874 3516 18880 3528
rect 18196 3488 18880 3516
rect 18196 3476 18202 3488
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 18969 3519 19027 3525
rect 18969 3485 18981 3519
rect 19015 3516 19027 3519
rect 19334 3516 19340 3528
rect 19015 3488 19340 3516
rect 19015 3485 19027 3488
rect 18969 3479 19027 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19610 3476 19616 3528
rect 19668 3476 19674 3528
rect 13688 3420 15240 3448
rect 13688 3408 13694 3420
rect 10321 3383 10379 3389
rect 10321 3380 10333 3383
rect 7852 3352 10333 3380
rect 10321 3349 10333 3352
rect 10367 3349 10379 3383
rect 10321 3343 10379 3349
rect 13078 3340 13084 3392
rect 13136 3380 13142 3392
rect 13998 3380 14004 3392
rect 13136 3352 14004 3380
rect 13136 3340 13142 3352
rect 13998 3340 14004 3352
rect 14056 3380 14062 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14056 3352 14933 3380
rect 14056 3340 14062 3352
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 15212 3380 15240 3420
rect 15473 3451 15531 3457
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 15519 3420 15884 3448
rect 17250 3420 17356 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 15746 3380 15752 3392
rect 15212 3352 15752 3380
rect 14921 3343 14979 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 15856 3380 15884 3420
rect 16482 3380 16488 3392
rect 15856 3352 16488 3380
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 17328 3380 17356 3420
rect 20438 3408 20444 3460
rect 20496 3408 20502 3460
rect 21910 3408 21916 3460
rect 21968 3408 21974 3460
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 17328 3352 17877 3380
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 17865 3343 17923 3349
rect 18138 3340 18144 3392
rect 18196 3340 18202 3392
rect 19886 3340 19892 3392
rect 19944 3380 19950 3392
rect 23308 3380 23336 3556
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3516 23443 3519
rect 23566 3516 23572 3528
rect 23431 3488 23572 3516
rect 23431 3485 23443 3488
rect 23385 3479 23443 3485
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 19944 3352 23336 3380
rect 19944 3340 19950 3352
rect 1104 3290 26312 3312
rect 1104 3238 4761 3290
rect 4813 3238 4825 3290
rect 4877 3238 4889 3290
rect 4941 3238 4953 3290
rect 5005 3238 5017 3290
rect 5069 3238 11063 3290
rect 11115 3238 11127 3290
rect 11179 3238 11191 3290
rect 11243 3238 11255 3290
rect 11307 3238 11319 3290
rect 11371 3238 17365 3290
rect 17417 3238 17429 3290
rect 17481 3238 17493 3290
rect 17545 3238 17557 3290
rect 17609 3238 17621 3290
rect 17673 3238 23667 3290
rect 23719 3238 23731 3290
rect 23783 3238 23795 3290
rect 23847 3238 23859 3290
rect 23911 3238 23923 3290
rect 23975 3238 26312 3290
rect 1104 3216 26312 3238
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6089 3179 6147 3185
rect 6089 3176 6101 3179
rect 5868 3148 6101 3176
rect 5868 3136 5874 3148
rect 6089 3145 6101 3148
rect 6135 3145 6147 3179
rect 6089 3139 6147 3145
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 6788 3148 6837 3176
rect 6788 3136 6794 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 8481 3179 8539 3185
rect 8481 3145 8493 3179
rect 8527 3176 8539 3179
rect 8754 3176 8760 3188
rect 8527 3148 8760 3176
rect 8527 3145 8539 3148
rect 8481 3139 8539 3145
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 11606 3176 11612 3188
rect 11379 3148 11612 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 14507 3179 14565 3185
rect 14507 3145 14519 3179
rect 14553 3176 14565 3179
rect 15194 3176 15200 3188
rect 14553 3148 15200 3176
rect 14553 3145 14565 3148
rect 14507 3139 14565 3145
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16393 3179 16451 3185
rect 16393 3145 16405 3179
rect 16439 3176 16451 3179
rect 17862 3176 17868 3188
rect 16439 3148 17868 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 20254 3136 20260 3188
rect 20312 3136 20318 3188
rect 20438 3136 20444 3188
rect 20496 3136 20502 3188
rect 21361 3179 21419 3185
rect 21361 3145 21373 3179
rect 21407 3176 21419 3179
rect 21910 3176 21916 3188
rect 21407 3148 21916 3176
rect 21407 3145 21419 3148
rect 21361 3139 21419 3145
rect 21910 3136 21916 3148
rect 21968 3136 21974 3188
rect 5626 3108 5632 3120
rect 4724 3080 5632 3108
rect 4724 3049 4752 3080
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 6362 3068 6368 3120
rect 6420 3068 6426 3120
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 10198 3111 10256 3117
rect 10198 3108 10210 3111
rect 10100 3080 10210 3108
rect 10100 3068 10106 3080
rect 10198 3077 10210 3080
rect 10244 3077 10256 3111
rect 10198 3071 10256 3077
rect 13814 3068 13820 3120
rect 13872 3068 13878 3120
rect 18138 3108 18144 3120
rect 18078 3080 18144 3108
rect 18138 3068 18144 3080
rect 18196 3068 18202 3120
rect 18509 3111 18567 3117
rect 18509 3077 18521 3111
rect 18555 3108 18567 3111
rect 18598 3108 18604 3120
rect 18555 3080 18604 3108
rect 18555 3077 18567 3080
rect 18509 3071 18567 3077
rect 18598 3068 18604 3080
rect 18656 3068 18662 3120
rect 20806 3108 20812 3120
rect 19996 3080 20812 3108
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4965 3043 5023 3049
rect 4965 3040 4977 3043
rect 4709 3003 4767 3009
rect 4816 3012 4977 3040
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 4816 2972 4844 3012
rect 4965 3009 4977 3012
rect 5011 3009 5023 3043
rect 4965 3003 5023 3009
rect 8662 3000 8668 3052
rect 8720 3000 8726 3052
rect 9950 3000 9956 3052
rect 10008 3000 10014 3052
rect 13078 3000 13084 3052
rect 13136 3000 13142 3052
rect 16298 3000 16304 3052
rect 16356 3000 16362 3052
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 19429 3043 19487 3049
rect 16715 3012 17172 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 4672 2944 4844 2972
rect 12713 2975 12771 2981
rect 4672 2932 4678 2944
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 12894 2972 12900 2984
rect 12759 2944 12900 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 17034 2932 17040 2984
rect 17092 2932 17098 2984
rect 17144 2972 17172 3012
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 19886 3040 19892 3052
rect 19475 3012 19892 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 19996 3049 20024 3080
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 19981 3003 20039 3009
rect 20088 3012 20361 3040
rect 17770 2972 17776 2984
rect 17144 2944 17776 2972
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 18874 2932 18880 2984
rect 18932 2972 18938 2984
rect 19705 2975 19763 2981
rect 19705 2972 19717 2975
rect 18932 2944 19717 2972
rect 18932 2932 18938 2944
rect 19705 2941 19717 2944
rect 19751 2972 19763 2975
rect 20088 2972 20116 3012
rect 20349 3009 20361 3012
rect 20395 3040 20407 3043
rect 21174 3040 21180 3052
rect 20395 3012 21180 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 21174 3000 21180 3012
rect 21232 3040 21238 3052
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 21232 3012 21281 3040
rect 21232 3000 21238 3012
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 19751 2944 20116 2972
rect 19751 2941 19763 2944
rect 19705 2935 19763 2941
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 20220 2944 20269 2972
rect 20220 2932 20226 2944
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 20257 2935 20315 2941
rect 6638 2864 6644 2916
rect 6696 2864 6702 2916
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 20073 2907 20131 2913
rect 20073 2904 20085 2907
rect 19484 2876 20085 2904
rect 19484 2864 19490 2876
rect 20073 2873 20085 2876
rect 20119 2873 20131 2907
rect 20073 2867 20131 2873
rect 1104 2746 26312 2768
rect 1104 2694 4101 2746
rect 4153 2694 4165 2746
rect 4217 2694 4229 2746
rect 4281 2694 4293 2746
rect 4345 2694 4357 2746
rect 4409 2694 10403 2746
rect 10455 2694 10467 2746
rect 10519 2694 10531 2746
rect 10583 2694 10595 2746
rect 10647 2694 10659 2746
rect 10711 2694 16705 2746
rect 16757 2694 16769 2746
rect 16821 2694 16833 2746
rect 16885 2694 16897 2746
rect 16949 2694 16961 2746
rect 17013 2694 23007 2746
rect 23059 2694 23071 2746
rect 23123 2694 23135 2746
rect 23187 2694 23199 2746
rect 23251 2694 23263 2746
rect 23315 2694 26312 2746
rect 1104 2672 26312 2694
rect 5994 2592 6000 2644
rect 6052 2592 6058 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 9122 2632 9128 2644
rect 8067 2604 9128 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 12066 2632 12072 2644
rect 11931 2604 12072 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 13814 2592 13820 2644
rect 13872 2592 13878 2644
rect 15565 2635 15623 2641
rect 15565 2601 15577 2635
rect 15611 2632 15623 2635
rect 16298 2632 16304 2644
rect 15611 2604 16304 2632
rect 15611 2601 15623 2604
rect 15565 2595 15623 2601
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 23566 2592 23572 2644
rect 23624 2632 23630 2644
rect 23937 2635 23995 2641
rect 23937 2632 23949 2635
rect 23624 2604 23949 2632
rect 23624 2592 23630 2604
rect 23937 2601 23949 2604
rect 23983 2601 23995 2635
rect 23937 2595 23995 2601
rect 17126 2564 17132 2576
rect 13740 2536 17132 2564
rect 11422 2496 11428 2508
rect 1504 2468 11428 2496
rect 1504 2437 1532 2468
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 1489 2431 1547 2437
rect 1489 2397 1501 2431
rect 1535 2397 1547 2431
rect 1489 2391 1547 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7800 2400 7849 2428
rect 7800 2388 7806 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 13740 2437 13768 2536
rect 17126 2524 17132 2536
rect 17184 2524 17190 2576
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14516 2468 20208 2496
rect 14516 2456 14522 2468
rect 13725 2431 13783 2437
rect 13725 2428 13737 2431
rect 12860 2400 13737 2428
rect 12860 2388 12866 2400
rect 13725 2397 13737 2400
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 20180 2437 20208 2468
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15528 2400 15761 2428
rect 15528 2388 15534 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2397 20223 2431
rect 20165 2391 20223 2397
rect 24026 2388 24032 2440
rect 24084 2428 24090 2440
rect 24121 2431 24179 2437
rect 24121 2428 24133 2431
rect 24084 2400 24133 2428
rect 24084 2388 24090 2400
rect 24121 2397 24133 2400
rect 24167 2397 24179 2431
rect 24121 2391 24179 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 72 2332 1869 2360
rect 72 2320 78 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 13446 2320 13452 2372
rect 13504 2360 13510 2372
rect 25593 2363 25651 2369
rect 25593 2360 25605 2363
rect 13504 2332 25605 2360
rect 13504 2320 13510 2332
rect 25593 2329 25605 2332
rect 25639 2329 25651 2363
rect 25593 2323 25651 2329
rect 4157 2295 4215 2301
rect 4157 2261 4169 2295
rect 4203 2292 4215 2295
rect 10870 2292 10876 2304
rect 4203 2264 10876 2292
rect 4203 2261 4215 2264
rect 4157 2255 4215 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 20036 2264 20269 2292
rect 20036 2252 20042 2264
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 24762 2252 24768 2304
rect 24820 2292 24826 2304
rect 25685 2295 25743 2301
rect 25685 2292 25697 2295
rect 24820 2264 25697 2292
rect 24820 2252 24826 2264
rect 25685 2261 25697 2264
rect 25731 2261 25743 2295
rect 25685 2255 25743 2261
rect 1104 2202 26312 2224
rect 1104 2150 4761 2202
rect 4813 2150 4825 2202
rect 4877 2150 4889 2202
rect 4941 2150 4953 2202
rect 5005 2150 5017 2202
rect 5069 2150 11063 2202
rect 11115 2150 11127 2202
rect 11179 2150 11191 2202
rect 11243 2150 11255 2202
rect 11307 2150 11319 2202
rect 11371 2150 17365 2202
rect 17417 2150 17429 2202
rect 17481 2150 17493 2202
rect 17545 2150 17557 2202
rect 17609 2150 17621 2202
rect 17673 2150 23667 2202
rect 23719 2150 23731 2202
rect 23783 2150 23795 2202
rect 23847 2150 23859 2202
rect 23911 2150 23923 2202
rect 23975 2150 26312 2202
rect 1104 2128 26312 2150
<< via1 >>
rect 4761 27174 4813 27226
rect 4825 27174 4877 27226
rect 4889 27174 4941 27226
rect 4953 27174 5005 27226
rect 5017 27174 5069 27226
rect 11063 27174 11115 27226
rect 11127 27174 11179 27226
rect 11191 27174 11243 27226
rect 11255 27174 11307 27226
rect 11319 27174 11371 27226
rect 17365 27174 17417 27226
rect 17429 27174 17481 27226
rect 17493 27174 17545 27226
rect 17557 27174 17609 27226
rect 17621 27174 17673 27226
rect 23667 27174 23719 27226
rect 23731 27174 23783 27226
rect 23795 27174 23847 27226
rect 23859 27174 23911 27226
rect 23923 27174 23975 27226
rect 3240 27072 3292 27124
rect 7104 27072 7156 27124
rect 11612 27072 11664 27124
rect 19340 27072 19392 27124
rect 23480 27115 23532 27124
rect 23480 27081 23489 27115
rect 23489 27081 23523 27115
rect 23523 27081 23532 27115
rect 23480 27072 23532 27081
rect 10784 27004 10836 27056
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 11520 26936 11572 26988
rect 12348 26936 12400 26988
rect 15476 26936 15528 26988
rect 19340 26936 19392 26988
rect 23388 26979 23440 26988
rect 23388 26945 23397 26979
rect 23397 26945 23431 26979
rect 23431 26945 23440 26979
rect 23388 26936 23440 26945
rect 2596 26732 2648 26784
rect 16304 26732 16356 26784
rect 4101 26630 4153 26682
rect 4165 26630 4217 26682
rect 4229 26630 4281 26682
rect 4293 26630 4345 26682
rect 4357 26630 4409 26682
rect 10403 26630 10455 26682
rect 10467 26630 10519 26682
rect 10531 26630 10583 26682
rect 10595 26630 10647 26682
rect 10659 26630 10711 26682
rect 16705 26630 16757 26682
rect 16769 26630 16821 26682
rect 16833 26630 16885 26682
rect 16897 26630 16949 26682
rect 16961 26630 17013 26682
rect 23007 26630 23059 26682
rect 23071 26630 23123 26682
rect 23135 26630 23187 26682
rect 23199 26630 23251 26682
rect 23263 26630 23315 26682
rect 9680 26503 9732 26512
rect 9680 26469 9689 26503
rect 9689 26469 9723 26503
rect 9723 26469 9732 26503
rect 9680 26460 9732 26469
rect 9864 26392 9916 26444
rect 13728 26392 13780 26444
rect 6552 26367 6604 26376
rect 6552 26333 6561 26367
rect 6561 26333 6595 26367
rect 6595 26333 6604 26367
rect 6552 26324 6604 26333
rect 8944 26324 8996 26376
rect 7472 26256 7524 26308
rect 9220 26299 9272 26308
rect 9220 26265 9229 26299
rect 9229 26265 9263 26299
rect 9263 26265 9272 26299
rect 9220 26256 9272 26265
rect 9404 26299 9456 26308
rect 9404 26265 9413 26299
rect 9413 26265 9447 26299
rect 9447 26265 9456 26299
rect 9404 26256 9456 26265
rect 9956 26367 10008 26376
rect 9956 26333 9965 26367
rect 9965 26333 9999 26367
rect 9999 26333 10008 26367
rect 9956 26324 10008 26333
rect 11888 26324 11940 26376
rect 12440 26367 12492 26376
rect 12440 26333 12449 26367
rect 12449 26333 12483 26367
rect 12483 26333 12492 26367
rect 12440 26324 12492 26333
rect 13820 26324 13872 26376
rect 18420 26392 18472 26444
rect 20720 26392 20772 26444
rect 15936 26324 15988 26376
rect 16580 26324 16632 26376
rect 8300 26231 8352 26240
rect 8300 26197 8309 26231
rect 8309 26197 8343 26231
rect 8343 26197 8352 26231
rect 8300 26188 8352 26197
rect 9588 26231 9640 26240
rect 9588 26197 9597 26231
rect 9597 26197 9631 26231
rect 9631 26197 9640 26231
rect 9588 26188 9640 26197
rect 10600 26256 10652 26308
rect 15476 26256 15528 26308
rect 17408 26367 17460 26376
rect 17408 26333 17417 26367
rect 17417 26333 17451 26367
rect 17451 26333 17460 26367
rect 17408 26324 17460 26333
rect 17776 26324 17828 26376
rect 19064 26324 19116 26376
rect 9772 26188 9824 26240
rect 10876 26188 10928 26240
rect 14648 26188 14700 26240
rect 17224 26188 17276 26240
rect 17408 26188 17460 26240
rect 20812 26256 20864 26308
rect 18788 26188 18840 26240
rect 4761 26086 4813 26138
rect 4825 26086 4877 26138
rect 4889 26086 4941 26138
rect 4953 26086 5005 26138
rect 5017 26086 5069 26138
rect 11063 26086 11115 26138
rect 11127 26086 11179 26138
rect 11191 26086 11243 26138
rect 11255 26086 11307 26138
rect 11319 26086 11371 26138
rect 17365 26086 17417 26138
rect 17429 26086 17481 26138
rect 17493 26086 17545 26138
rect 17557 26086 17609 26138
rect 17621 26086 17673 26138
rect 23667 26086 23719 26138
rect 23731 26086 23783 26138
rect 23795 26086 23847 26138
rect 23859 26086 23911 26138
rect 23923 26086 23975 26138
rect 6552 25916 6604 25968
rect 6920 25916 6972 25968
rect 8944 25916 8996 25968
rect 9128 25891 9180 25900
rect 9128 25857 9137 25891
rect 9137 25857 9171 25891
rect 9171 25857 9180 25891
rect 9128 25848 9180 25857
rect 9588 25916 9640 25968
rect 8760 25823 8812 25832
rect 8760 25789 8769 25823
rect 8769 25789 8803 25823
rect 8803 25789 8812 25823
rect 8760 25780 8812 25789
rect 9220 25780 9272 25832
rect 9588 25780 9640 25832
rect 9220 25644 9272 25696
rect 9404 25644 9456 25696
rect 10600 25891 10652 25900
rect 10600 25857 10609 25891
rect 10609 25857 10643 25891
rect 10643 25857 10652 25891
rect 10600 25848 10652 25857
rect 12808 25984 12860 26036
rect 13820 26027 13872 26036
rect 13820 25993 13829 26027
rect 13829 25993 13863 26027
rect 13863 25993 13872 26027
rect 13820 25984 13872 25993
rect 14648 25984 14700 26036
rect 15936 25984 15988 26036
rect 12716 25916 12768 25968
rect 15476 25916 15528 25968
rect 11888 25848 11940 25900
rect 10232 25644 10284 25696
rect 11612 25687 11664 25696
rect 11612 25653 11621 25687
rect 11621 25653 11655 25687
rect 11655 25653 11664 25687
rect 11612 25644 11664 25653
rect 13728 25891 13780 25900
rect 13728 25857 13737 25891
rect 13737 25857 13771 25891
rect 13771 25857 13780 25891
rect 13728 25848 13780 25857
rect 16304 25891 16356 25900
rect 16304 25857 16313 25891
rect 16313 25857 16347 25891
rect 16347 25857 16356 25891
rect 16304 25848 16356 25857
rect 18696 25984 18748 26036
rect 23388 25984 23440 26036
rect 20812 25916 20864 25968
rect 23572 25916 23624 25968
rect 17132 25848 17184 25900
rect 19432 25848 19484 25900
rect 15476 25780 15528 25832
rect 17040 25823 17092 25832
rect 17040 25789 17049 25823
rect 17049 25789 17083 25823
rect 17083 25789 17092 25823
rect 17040 25780 17092 25789
rect 19064 25780 19116 25832
rect 20076 25823 20128 25832
rect 20076 25789 20085 25823
rect 20085 25789 20119 25823
rect 20119 25789 20128 25823
rect 20076 25780 20128 25789
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22100 25848 22152 25857
rect 22652 25848 22704 25900
rect 22560 25823 22612 25832
rect 22560 25789 22569 25823
rect 22569 25789 22603 25823
rect 22603 25789 22612 25823
rect 22560 25780 22612 25789
rect 15844 25712 15896 25764
rect 13452 25644 13504 25696
rect 14004 25644 14056 25696
rect 16304 25644 16356 25696
rect 18236 25644 18288 25696
rect 18788 25687 18840 25696
rect 18788 25653 18797 25687
rect 18797 25653 18831 25687
rect 18831 25653 18840 25687
rect 18788 25644 18840 25653
rect 21272 25644 21324 25696
rect 24400 25644 24452 25696
rect 4101 25542 4153 25594
rect 4165 25542 4217 25594
rect 4229 25542 4281 25594
rect 4293 25542 4345 25594
rect 4357 25542 4409 25594
rect 10403 25542 10455 25594
rect 10467 25542 10519 25594
rect 10531 25542 10583 25594
rect 10595 25542 10647 25594
rect 10659 25542 10711 25594
rect 16705 25542 16757 25594
rect 16769 25542 16821 25594
rect 16833 25542 16885 25594
rect 16897 25542 16949 25594
rect 16961 25542 17013 25594
rect 23007 25542 23059 25594
rect 23071 25542 23123 25594
rect 23135 25542 23187 25594
rect 23199 25542 23251 25594
rect 23263 25542 23315 25594
rect 6920 25483 6972 25492
rect 6920 25449 6929 25483
rect 6929 25449 6963 25483
rect 6963 25449 6972 25483
rect 6920 25440 6972 25449
rect 7472 25483 7524 25492
rect 7472 25449 7481 25483
rect 7481 25449 7515 25483
rect 7515 25449 7524 25483
rect 7472 25440 7524 25449
rect 9036 25440 9088 25492
rect 9956 25440 10008 25492
rect 12716 25483 12768 25492
rect 12716 25449 12725 25483
rect 12725 25449 12759 25483
rect 12759 25449 12768 25483
rect 12716 25440 12768 25449
rect 12808 25440 12860 25492
rect 13728 25440 13780 25492
rect 15476 25483 15528 25492
rect 15476 25449 15485 25483
rect 15485 25449 15519 25483
rect 15519 25449 15528 25483
rect 15476 25440 15528 25449
rect 6552 25304 6604 25356
rect 8300 25304 8352 25356
rect 9864 25415 9916 25424
rect 9864 25381 9873 25415
rect 9873 25381 9907 25415
rect 9907 25381 9916 25415
rect 9864 25372 9916 25381
rect 10232 25372 10284 25424
rect 12440 25372 12492 25424
rect 13084 25372 13136 25424
rect 13544 25415 13596 25424
rect 13544 25381 13553 25415
rect 13553 25381 13587 25415
rect 13587 25381 13596 25415
rect 13544 25372 13596 25381
rect 6828 25279 6880 25288
rect 6828 25245 6837 25279
rect 6837 25245 6871 25279
rect 6871 25245 6880 25279
rect 6828 25236 6880 25245
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 9772 25304 9824 25356
rect 9496 25236 9548 25288
rect 9588 25279 9640 25288
rect 9588 25245 9597 25279
rect 9597 25245 9631 25279
rect 9631 25245 9640 25279
rect 9588 25236 9640 25245
rect 9680 25236 9732 25288
rect 10876 25304 10928 25356
rect 6000 25168 6052 25220
rect 6736 25211 6788 25220
rect 6736 25177 6745 25211
rect 6745 25177 6779 25211
rect 6779 25177 6788 25211
rect 6736 25168 6788 25177
rect 8760 25168 8812 25220
rect 9404 25211 9456 25220
rect 9404 25177 9413 25211
rect 9413 25177 9447 25211
rect 9447 25177 9456 25211
rect 9404 25168 9456 25177
rect 9956 25168 10008 25220
rect 10232 25279 10284 25288
rect 10232 25245 10241 25279
rect 10241 25245 10275 25279
rect 10275 25245 10284 25279
rect 10232 25236 10284 25245
rect 11612 25236 11664 25288
rect 12808 25236 12860 25288
rect 14832 25304 14884 25356
rect 6460 25100 6512 25152
rect 6552 25100 6604 25152
rect 10232 25100 10284 25152
rect 13820 25279 13872 25288
rect 13820 25245 13829 25279
rect 13829 25245 13863 25279
rect 13863 25245 13872 25279
rect 13820 25236 13872 25245
rect 14648 25236 14700 25288
rect 14924 25279 14976 25288
rect 14924 25245 14933 25279
rect 14933 25245 14967 25279
rect 14967 25245 14976 25279
rect 14924 25236 14976 25245
rect 16396 25304 16448 25356
rect 17868 25440 17920 25492
rect 23572 25440 23624 25492
rect 20812 25372 20864 25424
rect 17040 25304 17092 25356
rect 19432 25347 19484 25356
rect 19432 25313 19441 25347
rect 19441 25313 19475 25347
rect 19475 25313 19484 25347
rect 19432 25304 19484 25313
rect 21364 25347 21416 25356
rect 21364 25313 21373 25347
rect 21373 25313 21407 25347
rect 21407 25313 21416 25347
rect 21364 25304 21416 25313
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 15292 25236 15344 25245
rect 15752 25279 15804 25288
rect 15752 25245 15761 25279
rect 15761 25245 15795 25279
rect 15795 25245 15804 25279
rect 15752 25236 15804 25245
rect 16028 25279 16080 25288
rect 16028 25245 16037 25279
rect 16037 25245 16071 25279
rect 16071 25245 16080 25279
rect 16028 25236 16080 25245
rect 16948 25236 17000 25288
rect 17224 25236 17276 25288
rect 21272 25236 21324 25288
rect 22008 25236 22060 25288
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 14372 25100 14424 25152
rect 15016 25168 15068 25220
rect 19156 25168 19208 25220
rect 19708 25211 19760 25220
rect 19708 25177 19717 25211
rect 19717 25177 19751 25211
rect 19751 25177 19760 25211
rect 19708 25168 19760 25177
rect 20720 25168 20772 25220
rect 21364 25168 21416 25220
rect 24308 25236 24360 25288
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 25780 25279 25832 25288
rect 25780 25245 25789 25279
rect 25789 25245 25823 25279
rect 25823 25245 25832 25279
rect 25780 25236 25832 25245
rect 14924 25100 14976 25152
rect 16764 25100 16816 25152
rect 17040 25143 17092 25152
rect 17040 25109 17049 25143
rect 17049 25109 17083 25143
rect 17083 25109 17092 25143
rect 17040 25100 17092 25109
rect 17224 25100 17276 25152
rect 18880 25100 18932 25152
rect 21180 25143 21232 25152
rect 21180 25109 21189 25143
rect 21189 25109 21223 25143
rect 21223 25109 21232 25143
rect 21180 25100 21232 25109
rect 21824 25143 21876 25152
rect 21824 25109 21833 25143
rect 21833 25109 21867 25143
rect 21867 25109 21876 25143
rect 21824 25100 21876 25109
rect 22100 25100 22152 25152
rect 22744 25100 22796 25152
rect 23480 25143 23532 25152
rect 23480 25109 23489 25143
rect 23489 25109 23523 25143
rect 23523 25109 23532 25143
rect 23480 25100 23532 25109
rect 25044 25143 25096 25152
rect 25044 25109 25053 25143
rect 25053 25109 25087 25143
rect 25087 25109 25096 25143
rect 25044 25100 25096 25109
rect 25228 25100 25280 25152
rect 4761 24998 4813 25050
rect 4825 24998 4877 25050
rect 4889 24998 4941 25050
rect 4953 24998 5005 25050
rect 5017 24998 5069 25050
rect 11063 24998 11115 25050
rect 11127 24998 11179 25050
rect 11191 24998 11243 25050
rect 11255 24998 11307 25050
rect 11319 24998 11371 25050
rect 17365 24998 17417 25050
rect 17429 24998 17481 25050
rect 17493 24998 17545 25050
rect 17557 24998 17609 25050
rect 17621 24998 17673 25050
rect 23667 24998 23719 25050
rect 23731 24998 23783 25050
rect 23795 24998 23847 25050
rect 23859 24998 23911 25050
rect 23923 24998 23975 25050
rect 8116 24896 8168 24948
rect 9404 24939 9456 24948
rect 9404 24905 9429 24939
rect 9429 24905 9456 24939
rect 9404 24896 9456 24905
rect 6828 24828 6880 24880
rect 6000 24760 6052 24812
rect 6736 24803 6788 24812
rect 6736 24769 6745 24803
rect 6745 24769 6779 24803
rect 6779 24769 6788 24803
rect 6736 24760 6788 24769
rect 7564 24803 7616 24812
rect 7564 24769 7573 24803
rect 7573 24769 7607 24803
rect 7607 24769 7616 24803
rect 7564 24760 7616 24769
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 7840 24803 7892 24812
rect 7840 24769 7849 24803
rect 7849 24769 7883 24803
rect 7883 24769 7892 24803
rect 7840 24760 7892 24769
rect 8024 24803 8076 24812
rect 8024 24769 8033 24803
rect 8033 24769 8067 24803
rect 8067 24769 8076 24803
rect 8024 24760 8076 24769
rect 8300 24692 8352 24744
rect 9036 24760 9088 24812
rect 13084 24939 13136 24948
rect 13084 24905 13093 24939
rect 13093 24905 13127 24939
rect 13127 24905 13136 24939
rect 13084 24896 13136 24905
rect 13820 24896 13872 24948
rect 13544 24828 13596 24880
rect 7288 24556 7340 24608
rect 7472 24667 7524 24676
rect 7472 24633 7481 24667
rect 7481 24633 7515 24667
rect 7515 24633 7524 24667
rect 7472 24624 7524 24633
rect 8024 24624 8076 24676
rect 9680 24735 9732 24744
rect 9680 24701 9689 24735
rect 9689 24701 9723 24735
rect 9723 24701 9732 24735
rect 9680 24692 9732 24701
rect 10140 24760 10192 24812
rect 13636 24803 13688 24812
rect 13636 24769 13645 24803
rect 13645 24769 13679 24803
rect 13679 24769 13688 24803
rect 13636 24760 13688 24769
rect 13912 24760 13964 24812
rect 14924 24896 14976 24948
rect 15292 24896 15344 24948
rect 15752 24896 15804 24948
rect 16580 24896 16632 24948
rect 17132 24896 17184 24948
rect 17224 24896 17276 24948
rect 14372 24871 14424 24880
rect 14372 24837 14381 24871
rect 14381 24837 14415 24871
rect 14415 24837 14424 24871
rect 14372 24828 14424 24837
rect 15016 24828 15068 24880
rect 14464 24803 14516 24812
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 14648 24760 14700 24812
rect 14832 24760 14884 24812
rect 15200 24760 15252 24812
rect 19708 24939 19760 24948
rect 19708 24905 19717 24939
rect 19717 24905 19751 24939
rect 19751 24905 19760 24939
rect 19708 24896 19760 24905
rect 20076 24896 20128 24948
rect 16580 24760 16632 24812
rect 15752 24692 15804 24744
rect 16396 24692 16448 24744
rect 16488 24692 16540 24744
rect 16764 24803 16816 24812
rect 16764 24769 16773 24803
rect 16773 24769 16807 24803
rect 16807 24769 16816 24803
rect 16764 24760 16816 24769
rect 17040 24760 17092 24812
rect 17132 24803 17184 24812
rect 17132 24769 17141 24803
rect 17141 24769 17175 24803
rect 17175 24769 17184 24803
rect 17132 24760 17184 24769
rect 17224 24803 17276 24812
rect 17224 24769 17233 24803
rect 17233 24769 17267 24803
rect 17267 24769 17276 24803
rect 17224 24760 17276 24769
rect 17316 24803 17368 24812
rect 17316 24769 17325 24803
rect 17325 24769 17359 24803
rect 17359 24769 17368 24803
rect 17316 24760 17368 24769
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18144 24760 18196 24812
rect 18236 24803 18288 24812
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 18788 24828 18840 24880
rect 18696 24803 18748 24812
rect 18696 24769 18705 24803
rect 18705 24769 18739 24803
rect 18739 24769 18748 24803
rect 18696 24760 18748 24769
rect 18880 24803 18932 24812
rect 18880 24769 18889 24803
rect 18889 24769 18923 24803
rect 18923 24769 18932 24803
rect 18880 24760 18932 24769
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 19156 24803 19208 24812
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 22192 24896 22244 24948
rect 22468 24896 22520 24948
rect 20720 24871 20772 24880
rect 20720 24837 20729 24871
rect 20729 24837 20763 24871
rect 20763 24837 20772 24871
rect 20720 24828 20772 24837
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 20628 24803 20680 24812
rect 20628 24769 20637 24803
rect 20637 24769 20671 24803
rect 20671 24769 20680 24803
rect 20628 24760 20680 24769
rect 20812 24803 20864 24812
rect 21824 24828 21876 24880
rect 20812 24769 20847 24803
rect 20847 24769 20864 24803
rect 20812 24760 20864 24769
rect 21180 24760 21232 24812
rect 8208 24599 8260 24608
rect 8208 24565 8217 24599
rect 8217 24565 8251 24599
rect 8251 24565 8260 24599
rect 8208 24556 8260 24565
rect 8484 24599 8536 24608
rect 8484 24565 8493 24599
rect 8493 24565 8527 24599
rect 8527 24565 8536 24599
rect 8484 24556 8536 24565
rect 8944 24556 8996 24608
rect 9220 24556 9272 24608
rect 10324 24624 10376 24676
rect 13452 24624 13504 24676
rect 14924 24624 14976 24676
rect 19892 24735 19944 24744
rect 19892 24701 19901 24735
rect 19901 24701 19935 24735
rect 19935 24701 19944 24735
rect 19892 24692 19944 24701
rect 20076 24735 20128 24744
rect 20076 24701 20085 24735
rect 20085 24701 20119 24735
rect 20119 24701 20128 24735
rect 20076 24692 20128 24701
rect 22100 24803 22152 24812
rect 22100 24769 22109 24803
rect 22109 24769 22143 24803
rect 22143 24769 22152 24803
rect 22100 24760 22152 24769
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 22468 24760 22520 24812
rect 9680 24556 9732 24608
rect 12440 24556 12492 24608
rect 16396 24556 16448 24608
rect 17500 24624 17552 24676
rect 17868 24624 17920 24676
rect 17316 24556 17368 24608
rect 20812 24556 20864 24608
rect 21272 24624 21324 24676
rect 21456 24667 21508 24676
rect 21456 24633 21465 24667
rect 21465 24633 21499 24667
rect 21499 24633 21508 24667
rect 21456 24624 21508 24633
rect 4101 24454 4153 24506
rect 4165 24454 4217 24506
rect 4229 24454 4281 24506
rect 4293 24454 4345 24506
rect 4357 24454 4409 24506
rect 10403 24454 10455 24506
rect 10467 24454 10519 24506
rect 10531 24454 10583 24506
rect 10595 24454 10647 24506
rect 10659 24454 10711 24506
rect 16705 24454 16757 24506
rect 16769 24454 16821 24506
rect 16833 24454 16885 24506
rect 16897 24454 16949 24506
rect 16961 24454 17013 24506
rect 23007 24454 23059 24506
rect 23071 24454 23123 24506
rect 23135 24454 23187 24506
rect 23199 24454 23251 24506
rect 23263 24454 23315 24506
rect 6460 24352 6512 24404
rect 8024 24352 8076 24404
rect 8576 24395 8628 24404
rect 8576 24361 8585 24395
rect 8585 24361 8619 24395
rect 8619 24361 8628 24395
rect 8576 24352 8628 24361
rect 9312 24352 9364 24404
rect 14648 24395 14700 24404
rect 14648 24361 14657 24395
rect 14657 24361 14691 24395
rect 14691 24361 14700 24395
rect 14648 24352 14700 24361
rect 14924 24352 14976 24404
rect 15200 24352 15252 24404
rect 6552 24216 6604 24268
rect 6000 24191 6052 24200
rect 6000 24157 6009 24191
rect 6009 24157 6043 24191
rect 6043 24157 6052 24191
rect 6000 24148 6052 24157
rect 8208 24284 8260 24336
rect 8852 24284 8904 24336
rect 9036 24216 9088 24268
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 6552 24080 6604 24132
rect 8852 24148 8904 24200
rect 9312 24148 9364 24200
rect 9404 24191 9456 24200
rect 9404 24157 9413 24191
rect 9413 24157 9447 24191
rect 9447 24157 9456 24191
rect 9404 24148 9456 24157
rect 14740 24284 14792 24336
rect 15752 24395 15804 24404
rect 15752 24361 15761 24395
rect 15761 24361 15795 24395
rect 15795 24361 15804 24395
rect 15752 24352 15804 24361
rect 16028 24352 16080 24404
rect 16396 24352 16448 24404
rect 16580 24352 16632 24404
rect 17960 24352 18012 24404
rect 10232 24259 10284 24268
rect 10232 24225 10241 24259
rect 10241 24225 10275 24259
rect 10275 24225 10284 24259
rect 10232 24216 10284 24225
rect 12440 24259 12492 24268
rect 12440 24225 12449 24259
rect 12449 24225 12483 24259
rect 12483 24225 12492 24259
rect 12440 24216 12492 24225
rect 13636 24216 13688 24268
rect 14648 24216 14700 24268
rect 15660 24216 15712 24268
rect 9864 24191 9916 24200
rect 9864 24157 9873 24191
rect 9873 24157 9907 24191
rect 9907 24157 9916 24191
rect 9864 24148 9916 24157
rect 11612 24148 11664 24200
rect 11888 24148 11940 24200
rect 13820 24148 13872 24200
rect 14004 24148 14056 24200
rect 14740 24191 14792 24200
rect 14740 24157 14749 24191
rect 14749 24157 14783 24191
rect 14783 24157 14792 24191
rect 14740 24148 14792 24157
rect 8392 24123 8444 24132
rect 8392 24089 8401 24123
rect 8401 24089 8435 24123
rect 8435 24089 8444 24123
rect 8392 24080 8444 24089
rect 8484 24080 8536 24132
rect 7656 24012 7708 24064
rect 7748 24012 7800 24064
rect 8300 24012 8352 24064
rect 9496 24012 9548 24064
rect 9956 24012 10008 24064
rect 12992 24080 13044 24132
rect 15292 24123 15344 24132
rect 15292 24089 15301 24123
rect 15301 24089 15335 24123
rect 15335 24089 15344 24123
rect 15292 24080 15344 24089
rect 15568 24191 15620 24200
rect 15568 24157 15577 24191
rect 15577 24157 15611 24191
rect 15611 24157 15620 24191
rect 15568 24148 15620 24157
rect 12072 24012 12124 24064
rect 15752 24080 15804 24132
rect 17040 24284 17092 24336
rect 17224 24284 17276 24336
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 20720 24352 20772 24404
rect 21180 24352 21232 24404
rect 22376 24352 22428 24404
rect 22560 24352 22612 24404
rect 23388 24352 23440 24404
rect 20536 24284 20588 24336
rect 23480 24284 23532 24336
rect 16488 24148 16540 24200
rect 17040 24148 17092 24200
rect 18144 24148 18196 24200
rect 18880 24148 18932 24200
rect 20076 24148 20128 24200
rect 20904 24216 20956 24268
rect 22192 24216 22244 24268
rect 21088 24148 21140 24200
rect 21364 24148 21416 24200
rect 22284 24148 22336 24200
rect 20720 24080 20772 24132
rect 20812 24080 20864 24132
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 23572 24148 23624 24200
rect 19892 24012 19944 24064
rect 21364 24012 21416 24064
rect 22928 24080 22980 24132
rect 24308 24148 24360 24200
rect 23756 24123 23808 24132
rect 23756 24089 23765 24123
rect 23765 24089 23799 24123
rect 23799 24089 23808 24123
rect 23756 24080 23808 24089
rect 25044 24080 25096 24132
rect 23480 24012 23532 24064
rect 24492 24055 24544 24064
rect 24492 24021 24501 24055
rect 24501 24021 24535 24055
rect 24535 24021 24544 24055
rect 24492 24012 24544 24021
rect 4761 23910 4813 23962
rect 4825 23910 4877 23962
rect 4889 23910 4941 23962
rect 4953 23910 5005 23962
rect 5017 23910 5069 23962
rect 11063 23910 11115 23962
rect 11127 23910 11179 23962
rect 11191 23910 11243 23962
rect 11255 23910 11307 23962
rect 11319 23910 11371 23962
rect 17365 23910 17417 23962
rect 17429 23910 17481 23962
rect 17493 23910 17545 23962
rect 17557 23910 17609 23962
rect 17621 23910 17673 23962
rect 23667 23910 23719 23962
rect 23731 23910 23783 23962
rect 23795 23910 23847 23962
rect 23859 23910 23911 23962
rect 23923 23910 23975 23962
rect 6552 23851 6604 23860
rect 6552 23817 6561 23851
rect 6561 23817 6595 23851
rect 6595 23817 6604 23851
rect 6552 23808 6604 23817
rect 3700 23740 3752 23792
rect 5172 23783 5224 23792
rect 5172 23749 5181 23783
rect 5181 23749 5215 23783
rect 5215 23749 5224 23783
rect 5172 23740 5224 23749
rect 6000 23740 6052 23792
rect 7748 23808 7800 23860
rect 8852 23808 8904 23860
rect 9404 23808 9456 23860
rect 11612 23851 11664 23860
rect 11612 23817 11621 23851
rect 11621 23817 11655 23851
rect 11655 23817 11664 23851
rect 11612 23808 11664 23817
rect 12992 23808 13044 23860
rect 13636 23808 13688 23860
rect 16580 23808 16632 23860
rect 20904 23851 20956 23860
rect 20904 23817 20913 23851
rect 20913 23817 20947 23851
rect 20947 23817 20956 23851
rect 20904 23808 20956 23817
rect 22560 23808 22612 23860
rect 22928 23851 22980 23860
rect 22928 23817 22937 23851
rect 22937 23817 22971 23851
rect 22971 23817 22980 23851
rect 22928 23808 22980 23817
rect 3700 23511 3752 23520
rect 3700 23477 3709 23511
rect 3709 23477 3743 23511
rect 3743 23477 3752 23511
rect 3700 23468 3752 23477
rect 6460 23715 6512 23724
rect 6460 23681 6469 23715
rect 6469 23681 6503 23715
rect 6503 23681 6512 23715
rect 6460 23672 6512 23681
rect 7840 23740 7892 23792
rect 7288 23715 7340 23724
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 8208 23740 8260 23792
rect 8484 23672 8536 23724
rect 5540 23579 5592 23588
rect 5540 23545 5549 23579
rect 5549 23545 5583 23579
rect 5583 23545 5592 23579
rect 5540 23536 5592 23545
rect 7564 23604 7616 23656
rect 9312 23740 9364 23792
rect 9588 23740 9640 23792
rect 10140 23740 10192 23792
rect 8944 23715 8996 23724
rect 8944 23681 8953 23715
rect 8953 23681 8987 23715
rect 8987 23681 8996 23715
rect 8944 23672 8996 23681
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 9496 23672 9548 23724
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 10324 23672 10376 23724
rect 7472 23536 7524 23588
rect 7656 23536 7708 23588
rect 5632 23468 5684 23520
rect 8392 23536 8444 23588
rect 9036 23604 9088 23656
rect 8760 23579 8812 23588
rect 8760 23545 8773 23579
rect 8773 23545 8807 23579
rect 8807 23545 8812 23579
rect 8760 23536 8812 23545
rect 9128 23536 9180 23588
rect 8208 23468 8260 23520
rect 9588 23647 9640 23656
rect 9588 23613 9597 23647
rect 9597 23613 9631 23647
rect 9631 23613 9640 23647
rect 9588 23604 9640 23613
rect 9496 23579 9548 23588
rect 9496 23545 9505 23579
rect 9505 23545 9539 23579
rect 9539 23545 9548 23579
rect 9496 23536 9548 23545
rect 10140 23536 10192 23588
rect 10692 23647 10744 23656
rect 10692 23613 10701 23647
rect 10701 23613 10735 23647
rect 10735 23613 10744 23647
rect 10692 23604 10744 23613
rect 10784 23647 10836 23656
rect 10784 23613 10793 23647
rect 10793 23613 10827 23647
rect 10827 23613 10836 23647
rect 10784 23604 10836 23613
rect 11060 23672 11112 23724
rect 12900 23672 12952 23724
rect 13728 23672 13780 23724
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 14280 23715 14332 23724
rect 14280 23681 14289 23715
rect 14289 23681 14323 23715
rect 14323 23681 14332 23715
rect 14280 23672 14332 23681
rect 14648 23672 14700 23724
rect 14924 23740 14976 23792
rect 15292 23740 15344 23792
rect 15568 23783 15620 23792
rect 15568 23749 15577 23783
rect 15577 23749 15611 23783
rect 15611 23749 15620 23783
rect 15568 23740 15620 23749
rect 16304 23740 16356 23792
rect 21180 23740 21232 23792
rect 21364 23740 21416 23792
rect 12072 23604 12124 23656
rect 13912 23647 13964 23656
rect 13912 23613 13921 23647
rect 13921 23613 13955 23647
rect 13955 23613 13964 23647
rect 13912 23604 13964 23613
rect 15660 23604 15712 23656
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 12808 23536 12860 23588
rect 14464 23536 14516 23588
rect 22284 23740 22336 23792
rect 24492 23740 24544 23792
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 22560 23672 22612 23681
rect 23480 23672 23532 23724
rect 22652 23604 22704 23656
rect 9956 23511 10008 23520
rect 9956 23477 9965 23511
rect 9965 23477 9999 23511
rect 9999 23477 10008 23511
rect 9956 23468 10008 23477
rect 10048 23468 10100 23520
rect 10692 23468 10744 23520
rect 11704 23468 11756 23520
rect 16488 23468 16540 23520
rect 17040 23468 17092 23520
rect 20444 23468 20496 23520
rect 20720 23468 20772 23520
rect 21272 23511 21324 23520
rect 21272 23477 21281 23511
rect 21281 23477 21315 23511
rect 21315 23477 21324 23511
rect 21272 23468 21324 23477
rect 22928 23468 22980 23520
rect 23388 23468 23440 23520
rect 23664 23468 23716 23520
rect 4101 23366 4153 23418
rect 4165 23366 4217 23418
rect 4229 23366 4281 23418
rect 4293 23366 4345 23418
rect 4357 23366 4409 23418
rect 10403 23366 10455 23418
rect 10467 23366 10519 23418
rect 10531 23366 10583 23418
rect 10595 23366 10647 23418
rect 10659 23366 10711 23418
rect 16705 23366 16757 23418
rect 16769 23366 16821 23418
rect 16833 23366 16885 23418
rect 16897 23366 16949 23418
rect 16961 23366 17013 23418
rect 23007 23366 23059 23418
rect 23071 23366 23123 23418
rect 23135 23366 23187 23418
rect 23199 23366 23251 23418
rect 23263 23366 23315 23418
rect 5632 23264 5684 23316
rect 9036 23264 9088 23316
rect 9772 23264 9824 23316
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 19616 23264 19668 23316
rect 20628 23264 20680 23316
rect 20720 23264 20772 23316
rect 20996 23264 21048 23316
rect 9956 23196 10008 23248
rect 18052 23196 18104 23248
rect 19800 23196 19852 23248
rect 9128 23128 9180 23180
rect 12992 23128 13044 23180
rect 17960 23128 18012 23180
rect 3608 23060 3660 23112
rect 6000 23060 6052 23112
rect 9588 23060 9640 23112
rect 10048 23060 10100 23112
rect 16396 23060 16448 23112
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 4068 23035 4120 23044
rect 4068 23001 4077 23035
rect 4077 23001 4111 23035
rect 4111 23001 4120 23035
rect 4068 22992 4120 23001
rect 15936 22992 15988 23044
rect 6276 22967 6328 22976
rect 6276 22933 6285 22967
rect 6285 22933 6319 22967
rect 6319 22933 6328 22967
rect 6276 22924 6328 22933
rect 11980 22924 12032 22976
rect 16212 22924 16264 22976
rect 17132 22967 17184 22976
rect 17132 22933 17141 22967
rect 17141 22933 17175 22967
rect 17175 22933 17184 22967
rect 17132 22924 17184 22933
rect 17868 22992 17920 23044
rect 18512 23060 18564 23112
rect 19708 23060 19760 23112
rect 20168 23103 20220 23112
rect 20168 23069 20177 23103
rect 20177 23069 20211 23103
rect 20211 23069 20220 23103
rect 20168 23060 20220 23069
rect 20260 23062 20312 23114
rect 20444 23103 20496 23112
rect 20444 23069 20453 23103
rect 20453 23069 20487 23103
rect 20487 23069 20496 23103
rect 20444 23060 20496 23069
rect 20720 23128 20772 23180
rect 20996 23128 21048 23180
rect 21364 23196 21416 23248
rect 21272 23171 21324 23180
rect 21272 23137 21281 23171
rect 21281 23137 21315 23171
rect 21315 23137 21324 23171
rect 21272 23128 21324 23137
rect 20812 23060 20864 23112
rect 21088 23103 21140 23112
rect 21088 23069 21097 23103
rect 21097 23069 21131 23103
rect 21131 23069 21140 23103
rect 21088 23060 21140 23069
rect 19248 22992 19300 23044
rect 19892 22992 19944 23044
rect 22560 23264 22612 23316
rect 23388 23264 23440 23316
rect 23572 23264 23624 23316
rect 22376 23196 22428 23248
rect 22560 22992 22612 23044
rect 23664 23060 23716 23112
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 24216 23060 24268 23112
rect 18236 22924 18288 22976
rect 18328 22924 18380 22976
rect 20904 22924 20956 22976
rect 21364 22924 21416 22976
rect 4761 22822 4813 22874
rect 4825 22822 4877 22874
rect 4889 22822 4941 22874
rect 4953 22822 5005 22874
rect 5017 22822 5069 22874
rect 11063 22822 11115 22874
rect 11127 22822 11179 22874
rect 11191 22822 11243 22874
rect 11255 22822 11307 22874
rect 11319 22822 11371 22874
rect 17365 22822 17417 22874
rect 17429 22822 17481 22874
rect 17493 22822 17545 22874
rect 17557 22822 17609 22874
rect 17621 22822 17673 22874
rect 23667 22822 23719 22874
rect 23731 22822 23783 22874
rect 23795 22822 23847 22874
rect 23859 22822 23911 22874
rect 23923 22822 23975 22874
rect 4068 22763 4120 22772
rect 4068 22729 4077 22763
rect 4077 22729 4111 22763
rect 4111 22729 4120 22763
rect 4068 22720 4120 22729
rect 6276 22720 6328 22772
rect 6000 22695 6052 22704
rect 6000 22661 6009 22695
rect 6009 22661 6043 22695
rect 6043 22661 6052 22695
rect 6000 22652 6052 22661
rect 9220 22652 9272 22704
rect 9404 22652 9456 22704
rect 9772 22695 9824 22704
rect 9772 22661 9797 22695
rect 9797 22661 9824 22695
rect 9956 22763 10008 22772
rect 9956 22729 9965 22763
rect 9965 22729 9999 22763
rect 9999 22729 10008 22763
rect 9956 22720 10008 22729
rect 10784 22720 10836 22772
rect 11704 22763 11756 22772
rect 11704 22729 11729 22763
rect 11729 22729 11756 22763
rect 11704 22720 11756 22729
rect 11980 22720 12032 22772
rect 12072 22720 12124 22772
rect 12992 22720 13044 22772
rect 9772 22652 9824 22661
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 6276 22584 6328 22636
rect 6460 22584 6512 22636
rect 11612 22584 11664 22636
rect 11980 22584 12032 22636
rect 6184 22448 6236 22500
rect 12532 22516 12584 22568
rect 15016 22584 15068 22636
rect 15660 22652 15712 22704
rect 16304 22652 16356 22704
rect 17040 22695 17092 22704
rect 17040 22661 17049 22695
rect 17049 22661 17083 22695
rect 17083 22661 17092 22695
rect 17040 22652 17092 22661
rect 12808 22559 12860 22568
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 12992 22516 13044 22568
rect 16396 22584 16448 22636
rect 18144 22720 18196 22772
rect 19708 22763 19760 22772
rect 19708 22729 19717 22763
rect 19717 22729 19751 22763
rect 19751 22729 19760 22763
rect 19708 22720 19760 22729
rect 20076 22720 20128 22772
rect 21456 22720 21508 22772
rect 22560 22763 22612 22772
rect 22560 22729 22569 22763
rect 22569 22729 22603 22763
rect 22603 22729 22612 22763
rect 22560 22720 22612 22729
rect 18604 22652 18656 22704
rect 17132 22516 17184 22568
rect 17316 22516 17368 22568
rect 18328 22584 18380 22636
rect 18512 22584 18564 22636
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 19800 22652 19852 22704
rect 21548 22652 21600 22704
rect 23756 22652 23808 22704
rect 24216 22652 24268 22704
rect 19708 22627 19760 22636
rect 19708 22593 19717 22627
rect 19717 22593 19751 22627
rect 19751 22593 19760 22627
rect 19708 22584 19760 22593
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 10324 22423 10376 22432
rect 10324 22389 10333 22423
rect 10333 22389 10367 22423
rect 10367 22389 10376 22423
rect 10324 22380 10376 22389
rect 10876 22380 10928 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 12440 22423 12492 22432
rect 12440 22389 12449 22423
rect 12449 22389 12483 22423
rect 12483 22389 12492 22423
rect 12440 22380 12492 22389
rect 12808 22380 12860 22432
rect 15200 22491 15252 22500
rect 15200 22457 15209 22491
rect 15209 22457 15243 22491
rect 15243 22457 15252 22491
rect 15200 22448 15252 22457
rect 16028 22448 16080 22500
rect 17776 22448 17828 22500
rect 18328 22448 18380 22500
rect 19616 22516 19668 22568
rect 20352 22516 20404 22568
rect 20996 22516 21048 22568
rect 22284 22516 22336 22568
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 22928 22584 22980 22636
rect 19432 22448 19484 22500
rect 21364 22448 21416 22500
rect 13728 22380 13780 22432
rect 15568 22423 15620 22432
rect 15568 22389 15577 22423
rect 15577 22389 15611 22423
rect 15611 22389 15620 22423
rect 15568 22380 15620 22389
rect 16120 22380 16172 22432
rect 16304 22380 16356 22432
rect 17040 22423 17092 22432
rect 17040 22389 17049 22423
rect 17049 22389 17083 22423
rect 17083 22389 17092 22423
rect 17040 22380 17092 22389
rect 17224 22423 17276 22432
rect 17224 22389 17233 22423
rect 17233 22389 17267 22423
rect 17267 22389 17276 22423
rect 17224 22380 17276 22389
rect 17684 22423 17736 22432
rect 17684 22389 17693 22423
rect 17693 22389 17727 22423
rect 17727 22389 17736 22423
rect 17684 22380 17736 22389
rect 18880 22423 18932 22432
rect 18880 22389 18889 22423
rect 18889 22389 18923 22423
rect 18923 22389 18932 22423
rect 18880 22380 18932 22389
rect 19708 22380 19760 22432
rect 21088 22380 21140 22432
rect 24032 22516 24084 22568
rect 4101 22278 4153 22330
rect 4165 22278 4217 22330
rect 4229 22278 4281 22330
rect 4293 22278 4345 22330
rect 4357 22278 4409 22330
rect 10403 22278 10455 22330
rect 10467 22278 10519 22330
rect 10531 22278 10583 22330
rect 10595 22278 10647 22330
rect 10659 22278 10711 22330
rect 16705 22278 16757 22330
rect 16769 22278 16821 22330
rect 16833 22278 16885 22330
rect 16897 22278 16949 22330
rect 16961 22278 17013 22330
rect 23007 22278 23059 22330
rect 23071 22278 23123 22330
rect 23135 22278 23187 22330
rect 23199 22278 23251 22330
rect 23263 22278 23315 22330
rect 11336 22176 11388 22228
rect 11980 22108 12032 22160
rect 15936 22219 15988 22228
rect 15936 22185 15945 22219
rect 15945 22185 15979 22219
rect 15979 22185 15988 22219
rect 15936 22176 15988 22185
rect 17132 22176 17184 22228
rect 17224 22176 17276 22228
rect 17868 22176 17920 22228
rect 17776 22108 17828 22160
rect 18328 22151 18380 22160
rect 18328 22117 18337 22151
rect 18337 22117 18371 22151
rect 18371 22117 18380 22151
rect 18328 22108 18380 22117
rect 18512 22219 18564 22228
rect 18512 22185 18521 22219
rect 18521 22185 18555 22219
rect 18555 22185 18564 22219
rect 18512 22176 18564 22185
rect 19248 22176 19300 22228
rect 20076 22176 20128 22228
rect 4160 21972 4212 22024
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 5908 22015 5960 22024
rect 5908 21981 5917 22015
rect 5917 21981 5951 22015
rect 5951 21981 5960 22015
rect 5908 21972 5960 21981
rect 6736 21972 6788 22024
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 9312 21972 9364 22024
rect 12716 22040 12768 22092
rect 12992 22040 13044 22092
rect 11980 21972 12032 22024
rect 12072 22015 12124 22024
rect 12072 21981 12081 22015
rect 12081 21981 12115 22015
rect 12115 21981 12124 22015
rect 12072 21972 12124 21981
rect 7472 21904 7524 21956
rect 3792 21836 3844 21888
rect 6644 21836 6696 21888
rect 7104 21836 7156 21888
rect 10324 21904 10376 21956
rect 13084 21904 13136 21956
rect 15016 22040 15068 22092
rect 16120 22040 16172 22092
rect 13912 21972 13964 22024
rect 14280 21972 14332 22024
rect 15292 21972 15344 22024
rect 16028 21904 16080 21956
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 16856 22015 16908 22024
rect 16856 21981 16865 22015
rect 16865 21981 16899 22015
rect 16899 21981 16908 22015
rect 16856 21972 16908 21981
rect 17316 22040 17368 22092
rect 19800 22083 19852 22092
rect 19800 22049 19809 22083
rect 19809 22049 19843 22083
rect 19843 22049 19852 22083
rect 19800 22040 19852 22049
rect 21548 22083 21600 22092
rect 21548 22049 21557 22083
rect 21557 22049 21591 22083
rect 21591 22049 21600 22083
rect 21548 22040 21600 22049
rect 23756 22083 23808 22092
rect 23756 22049 23765 22083
rect 23765 22049 23799 22083
rect 23799 22049 23808 22083
rect 23756 22040 23808 22049
rect 17776 22015 17828 22024
rect 17776 21981 17785 22015
rect 17785 21981 17819 22015
rect 17819 21981 17828 22015
rect 17776 21972 17828 21981
rect 19248 21972 19300 22024
rect 19524 21972 19576 22024
rect 24308 21972 24360 22024
rect 17868 21904 17920 21956
rect 18052 21904 18104 21956
rect 18604 21947 18656 21956
rect 18604 21913 18613 21947
rect 18613 21913 18647 21947
rect 18647 21913 18656 21947
rect 18604 21904 18656 21913
rect 8944 21879 8996 21888
rect 8944 21845 8953 21879
rect 8953 21845 8987 21879
rect 8987 21845 8996 21879
rect 8944 21836 8996 21845
rect 11612 21836 11664 21888
rect 12532 21836 12584 21888
rect 13636 21836 13688 21888
rect 14464 21836 14516 21888
rect 16212 21836 16264 21888
rect 16580 21836 16632 21888
rect 17040 21836 17092 21888
rect 18972 21879 19024 21888
rect 18972 21845 18981 21879
rect 18981 21845 19015 21879
rect 19015 21845 19024 21879
rect 18972 21836 19024 21845
rect 19708 21947 19760 21956
rect 19708 21913 19717 21947
rect 19717 21913 19751 21947
rect 19751 21913 19760 21947
rect 19708 21904 19760 21913
rect 21088 21836 21140 21888
rect 4761 21734 4813 21786
rect 4825 21734 4877 21786
rect 4889 21734 4941 21786
rect 4953 21734 5005 21786
rect 5017 21734 5069 21786
rect 11063 21734 11115 21786
rect 11127 21734 11179 21786
rect 11191 21734 11243 21786
rect 11255 21734 11307 21786
rect 11319 21734 11371 21786
rect 17365 21734 17417 21786
rect 17429 21734 17481 21786
rect 17493 21734 17545 21786
rect 17557 21734 17609 21786
rect 17621 21734 17673 21786
rect 23667 21734 23719 21786
rect 23731 21734 23783 21786
rect 23795 21734 23847 21786
rect 23859 21734 23911 21786
rect 23923 21734 23975 21786
rect 3608 21632 3660 21684
rect 5540 21632 5592 21684
rect 9128 21632 9180 21684
rect 2504 21564 2556 21616
rect 3516 21564 3568 21616
rect 6644 21607 6696 21616
rect 6644 21573 6653 21607
rect 6653 21573 6687 21607
rect 6687 21573 6696 21607
rect 6644 21564 6696 21573
rect 7104 21564 7156 21616
rect 8944 21564 8996 21616
rect 10876 21564 10928 21616
rect 12440 21632 12492 21684
rect 13728 21632 13780 21684
rect 16304 21632 16356 21684
rect 17132 21632 17184 21684
rect 14372 21564 14424 21616
rect 16120 21564 16172 21616
rect 18052 21564 18104 21616
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 8668 21496 8720 21548
rect 1400 21428 1452 21480
rect 2136 21428 2188 21480
rect 2872 21360 2924 21412
rect 3884 21471 3936 21480
rect 3884 21437 3893 21471
rect 3893 21437 3927 21471
rect 3927 21437 3936 21471
rect 3884 21428 3936 21437
rect 5172 21428 5224 21480
rect 5632 21428 5684 21480
rect 6368 21471 6420 21480
rect 6368 21437 6377 21471
rect 6377 21437 6411 21471
rect 6411 21437 6420 21471
rect 6368 21428 6420 21437
rect 3608 21292 3660 21344
rect 3976 21292 4028 21344
rect 8024 21360 8076 21412
rect 7656 21292 7708 21344
rect 12072 21496 12124 21548
rect 9312 21471 9364 21480
rect 9312 21437 9321 21471
rect 9321 21437 9355 21471
rect 9355 21437 9364 21471
rect 9312 21428 9364 21437
rect 14464 21496 14516 21548
rect 14740 21496 14792 21548
rect 15292 21539 15344 21548
rect 15292 21505 15301 21539
rect 15301 21505 15335 21539
rect 15335 21505 15344 21539
rect 15292 21496 15344 21505
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 18972 21564 19024 21616
rect 18236 21496 18288 21548
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 25780 21539 25832 21548
rect 25780 21505 25789 21539
rect 25789 21505 25823 21539
rect 25823 21505 25832 21539
rect 25780 21496 25832 21505
rect 14096 21428 14148 21480
rect 14280 21360 14332 21412
rect 16856 21428 16908 21480
rect 17500 21428 17552 21480
rect 19984 21428 20036 21480
rect 21364 21428 21416 21480
rect 15108 21360 15160 21412
rect 9772 21292 9824 21344
rect 13636 21292 13688 21344
rect 15568 21292 15620 21344
rect 16028 21292 16080 21344
rect 17868 21292 17920 21344
rect 18144 21360 18196 21412
rect 19800 21292 19852 21344
rect 25964 21335 26016 21344
rect 25964 21301 25973 21335
rect 25973 21301 26007 21335
rect 26007 21301 26016 21335
rect 25964 21292 26016 21301
rect 4101 21190 4153 21242
rect 4165 21190 4217 21242
rect 4229 21190 4281 21242
rect 4293 21190 4345 21242
rect 4357 21190 4409 21242
rect 10403 21190 10455 21242
rect 10467 21190 10519 21242
rect 10531 21190 10583 21242
rect 10595 21190 10647 21242
rect 10659 21190 10711 21242
rect 16705 21190 16757 21242
rect 16769 21190 16821 21242
rect 16833 21190 16885 21242
rect 16897 21190 16949 21242
rect 16961 21190 17013 21242
rect 23007 21190 23059 21242
rect 23071 21190 23123 21242
rect 23135 21190 23187 21242
rect 23199 21190 23251 21242
rect 23263 21190 23315 21242
rect 2136 21131 2188 21140
rect 2136 21097 2145 21131
rect 2145 21097 2179 21131
rect 2179 21097 2188 21131
rect 2136 21088 2188 21097
rect 2504 21131 2556 21140
rect 2504 21097 2513 21131
rect 2513 21097 2547 21131
rect 2547 21097 2556 21131
rect 2504 21088 2556 21097
rect 2780 21088 2832 21140
rect 3424 21088 3476 21140
rect 3516 21131 3568 21140
rect 3516 21097 3525 21131
rect 3525 21097 3559 21131
rect 3559 21097 3568 21131
rect 3516 21088 3568 21097
rect 3884 21088 3936 21140
rect 4344 21088 4396 21140
rect 5264 21088 5316 21140
rect 5632 21088 5684 21140
rect 5172 21020 5224 21072
rect 5908 21088 5960 21140
rect 6920 21088 6972 21140
rect 8024 21131 8076 21140
rect 8024 21097 8033 21131
rect 8033 21097 8067 21131
rect 8067 21097 8076 21131
rect 8024 21088 8076 21097
rect 8760 21088 8812 21140
rect 11888 21131 11940 21140
rect 11888 21097 11897 21131
rect 11897 21097 11931 21131
rect 11931 21097 11940 21131
rect 11888 21088 11940 21097
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 14372 21131 14424 21140
rect 14372 21097 14381 21131
rect 14381 21097 14415 21131
rect 14415 21097 14424 21131
rect 14372 21088 14424 21097
rect 17224 21088 17276 21140
rect 17960 21088 18012 21140
rect 18604 21088 18656 21140
rect 2872 20952 2924 21004
rect 3332 20952 3384 21004
rect 7288 21020 7340 21072
rect 7472 21020 7524 21072
rect 940 20884 992 20936
rect 2320 20884 2372 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 5540 20952 5592 21004
rect 6644 20952 6696 21004
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 5264 20884 5316 20936
rect 7656 20884 7708 20936
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 5816 20816 5868 20868
rect 5908 20859 5960 20868
rect 5908 20825 5917 20859
rect 5917 20825 5951 20859
rect 5951 20825 5960 20859
rect 5908 20816 5960 20825
rect 9404 20995 9456 21004
rect 9404 20961 9413 20995
rect 9413 20961 9447 20995
rect 9447 20961 9456 20995
rect 9404 20952 9456 20961
rect 14096 21020 14148 21072
rect 19708 21088 19760 21140
rect 21364 21131 21416 21140
rect 21364 21097 21373 21131
rect 21373 21097 21407 21131
rect 21407 21097 21416 21131
rect 21364 21088 21416 21097
rect 11612 20952 11664 21004
rect 15200 20952 15252 21004
rect 16120 20952 16172 21004
rect 5540 20791 5592 20800
rect 5540 20757 5549 20791
rect 5549 20757 5583 20791
rect 5583 20757 5592 20791
rect 5540 20748 5592 20757
rect 6736 20748 6788 20800
rect 8668 20884 8720 20936
rect 12900 20884 12952 20936
rect 13268 20884 13320 20936
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 10968 20816 11020 20868
rect 15844 20816 15896 20868
rect 16856 20952 16908 21004
rect 19616 20995 19668 21004
rect 19616 20961 19625 20995
rect 19625 20961 19659 20995
rect 19659 20961 19668 20995
rect 19616 20952 19668 20961
rect 16580 20884 16632 20936
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 18052 20884 18104 20936
rect 24032 20952 24084 21004
rect 17132 20816 17184 20868
rect 19892 20859 19944 20868
rect 19892 20825 19901 20859
rect 19901 20825 19935 20859
rect 19935 20825 19944 20859
rect 19892 20816 19944 20825
rect 23480 20884 23532 20936
rect 24308 20884 24360 20936
rect 24768 20884 24820 20936
rect 16580 20791 16632 20800
rect 16580 20757 16589 20791
rect 16589 20757 16623 20791
rect 16623 20757 16632 20791
rect 16580 20748 16632 20757
rect 23388 20791 23440 20800
rect 23388 20757 23397 20791
rect 23397 20757 23431 20791
rect 23431 20757 23440 20791
rect 23388 20748 23440 20757
rect 24032 20748 24084 20800
rect 4761 20646 4813 20698
rect 4825 20646 4877 20698
rect 4889 20646 4941 20698
rect 4953 20646 5005 20698
rect 5017 20646 5069 20698
rect 11063 20646 11115 20698
rect 11127 20646 11179 20698
rect 11191 20646 11243 20698
rect 11255 20646 11307 20698
rect 11319 20646 11371 20698
rect 17365 20646 17417 20698
rect 17429 20646 17481 20698
rect 17493 20646 17545 20698
rect 17557 20646 17609 20698
rect 17621 20646 17673 20698
rect 23667 20646 23719 20698
rect 23731 20646 23783 20698
rect 23795 20646 23847 20698
rect 23859 20646 23911 20698
rect 23923 20646 23975 20698
rect 3424 20587 3476 20596
rect 3424 20553 3433 20587
rect 3433 20553 3467 20587
rect 3467 20553 3476 20587
rect 3424 20544 3476 20553
rect 5264 20544 5316 20596
rect 6920 20544 6972 20596
rect 7472 20587 7524 20596
rect 7472 20553 7481 20587
rect 7481 20553 7515 20587
rect 7515 20553 7524 20587
rect 7472 20544 7524 20553
rect 2872 20408 2924 20460
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 5172 20519 5224 20528
rect 5172 20485 5181 20519
rect 5181 20485 5215 20519
rect 5215 20485 5224 20519
rect 5172 20476 5224 20485
rect 3516 20340 3568 20392
rect 4344 20408 4396 20460
rect 4804 20408 4856 20460
rect 6368 20476 6420 20528
rect 9312 20544 9364 20596
rect 10048 20544 10100 20596
rect 10784 20544 10836 20596
rect 19616 20544 19668 20596
rect 5540 20408 5592 20460
rect 6276 20408 6328 20460
rect 6552 20451 6604 20460
rect 6552 20417 6561 20451
rect 6561 20417 6595 20451
rect 6595 20417 6604 20451
rect 6552 20408 6604 20417
rect 9220 20476 9272 20528
rect 10140 20476 10192 20528
rect 10968 20476 11020 20528
rect 12440 20476 12492 20528
rect 17224 20476 17276 20528
rect 5448 20340 5500 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 6736 20383 6788 20392
rect 6736 20349 6745 20383
rect 6745 20349 6779 20383
rect 6779 20349 6788 20383
rect 6736 20340 6788 20349
rect 6828 20340 6880 20392
rect 11428 20408 11480 20460
rect 8484 20383 8536 20392
rect 8484 20349 8493 20383
rect 8493 20349 8527 20383
rect 8527 20349 8536 20383
rect 8484 20340 8536 20349
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 4436 20204 4488 20256
rect 4528 20204 4580 20256
rect 4712 20204 4764 20256
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 6092 20247 6144 20256
rect 6092 20213 6101 20247
rect 6101 20213 6135 20247
rect 6135 20213 6144 20247
rect 6092 20204 6144 20213
rect 6276 20204 6328 20256
rect 6736 20204 6788 20256
rect 9588 20272 9640 20324
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 13636 20451 13688 20460
rect 13636 20417 13645 20451
rect 13645 20417 13679 20451
rect 13679 20417 13688 20451
rect 13636 20408 13688 20417
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 22008 20476 22060 20528
rect 17960 20451 18012 20460
rect 17960 20417 17969 20451
rect 17969 20417 18003 20451
rect 18003 20417 18012 20451
rect 17960 20408 18012 20417
rect 19064 20408 19116 20460
rect 20444 20408 20496 20460
rect 21456 20408 21508 20460
rect 24032 20476 24084 20528
rect 24768 20519 24820 20528
rect 24768 20485 24777 20519
rect 24777 20485 24811 20519
rect 24811 20485 24820 20519
rect 24768 20476 24820 20485
rect 23388 20408 23440 20460
rect 13268 20272 13320 20324
rect 17776 20340 17828 20392
rect 20628 20383 20680 20392
rect 20628 20349 20637 20383
rect 20637 20349 20671 20383
rect 20671 20349 20680 20383
rect 20628 20340 20680 20349
rect 20904 20340 20956 20392
rect 21640 20340 21692 20392
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 15936 20204 15988 20256
rect 16028 20247 16080 20256
rect 16028 20213 16037 20247
rect 16037 20213 16071 20247
rect 16071 20213 16080 20247
rect 16028 20204 16080 20213
rect 16304 20204 16356 20256
rect 16580 20204 16632 20256
rect 18052 20247 18104 20256
rect 18052 20213 18061 20247
rect 18061 20213 18095 20247
rect 18095 20213 18104 20247
rect 18052 20204 18104 20213
rect 18236 20272 18288 20324
rect 25136 20340 25188 20392
rect 18512 20204 18564 20256
rect 20996 20204 21048 20256
rect 21272 20247 21324 20256
rect 21272 20213 21281 20247
rect 21281 20213 21315 20247
rect 21315 20213 21324 20247
rect 21272 20204 21324 20213
rect 21364 20204 21416 20256
rect 4101 20102 4153 20154
rect 4165 20102 4217 20154
rect 4229 20102 4281 20154
rect 4293 20102 4345 20154
rect 4357 20102 4409 20154
rect 10403 20102 10455 20154
rect 10467 20102 10519 20154
rect 10531 20102 10583 20154
rect 10595 20102 10647 20154
rect 10659 20102 10711 20154
rect 16705 20102 16757 20154
rect 16769 20102 16821 20154
rect 16833 20102 16885 20154
rect 16897 20102 16949 20154
rect 16961 20102 17013 20154
rect 23007 20102 23059 20154
rect 23071 20102 23123 20154
rect 23135 20102 23187 20154
rect 23199 20102 23251 20154
rect 23263 20102 23315 20154
rect 2872 20000 2924 20052
rect 3424 20000 3476 20052
rect 4436 20000 4488 20052
rect 4804 20000 4856 20052
rect 5356 20000 5408 20052
rect 5724 20043 5776 20052
rect 5724 20009 5733 20043
rect 5733 20009 5767 20043
rect 5767 20009 5776 20043
rect 5724 20000 5776 20009
rect 5908 20043 5960 20052
rect 5908 20009 5917 20043
rect 5917 20009 5951 20043
rect 5951 20009 5960 20043
rect 5908 20000 5960 20009
rect 6920 20000 6972 20052
rect 9220 20043 9272 20052
rect 9220 20009 9229 20043
rect 9229 20009 9263 20043
rect 9263 20009 9272 20043
rect 9220 20000 9272 20009
rect 6368 19932 6420 19984
rect 6644 19932 6696 19984
rect 9956 20000 10008 20052
rect 11428 20043 11480 20052
rect 11428 20009 11437 20043
rect 11437 20009 11471 20043
rect 11471 20009 11480 20043
rect 11428 20000 11480 20009
rect 11704 20000 11756 20052
rect 12348 20000 12400 20052
rect 1676 19660 1728 19712
rect 3516 19864 3568 19916
rect 5172 19907 5224 19916
rect 5172 19873 5181 19907
rect 5181 19873 5215 19907
rect 5215 19873 5224 19907
rect 5172 19864 5224 19873
rect 5448 19864 5500 19916
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 2780 19796 2832 19805
rect 2964 19839 3016 19848
rect 2964 19805 2973 19839
rect 2973 19805 3007 19839
rect 3007 19805 3016 19839
rect 2964 19796 3016 19805
rect 3332 19839 3384 19848
rect 3332 19805 3341 19839
rect 3341 19805 3375 19839
rect 3375 19805 3384 19839
rect 3332 19796 3384 19805
rect 3424 19839 3476 19848
rect 3424 19805 3433 19839
rect 3433 19805 3467 19839
rect 3467 19805 3476 19839
rect 3424 19796 3476 19805
rect 4712 19796 4764 19848
rect 5724 19796 5776 19848
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 7104 19864 7156 19916
rect 7656 19864 7708 19916
rect 7288 19839 7340 19848
rect 7288 19805 7297 19839
rect 7297 19805 7331 19839
rect 7331 19805 7340 19839
rect 7288 19796 7340 19805
rect 12624 19932 12676 19984
rect 9312 19864 9364 19916
rect 13636 19864 13688 19916
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 9588 19796 9640 19805
rect 11428 19796 11480 19848
rect 4436 19660 4488 19712
rect 4528 19660 4580 19712
rect 6644 19728 6696 19780
rect 7932 19728 7984 19780
rect 5356 19660 5408 19712
rect 6000 19660 6052 19712
rect 6736 19660 6788 19712
rect 8024 19703 8076 19712
rect 8024 19669 8033 19703
rect 8033 19669 8067 19703
rect 8067 19669 8076 19703
rect 8024 19660 8076 19669
rect 12716 19796 12768 19848
rect 13452 19796 13504 19848
rect 14004 19728 14056 19780
rect 16488 19932 16540 19984
rect 16580 19932 16632 19984
rect 19892 20000 19944 20052
rect 25964 20000 26016 20052
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 18236 19796 18288 19848
rect 19156 19796 19208 19848
rect 20168 19796 20220 19848
rect 21824 19932 21876 19984
rect 20444 19907 20496 19916
rect 20444 19873 20453 19907
rect 20453 19873 20487 19907
rect 20487 19873 20496 19907
rect 20444 19864 20496 19873
rect 20996 19864 21048 19916
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22008 19864 22060 19873
rect 22284 19864 22336 19916
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 20444 19728 20496 19780
rect 21272 19839 21324 19848
rect 21272 19805 21281 19839
rect 21281 19805 21315 19839
rect 21315 19805 21324 19839
rect 21272 19796 21324 19805
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 21180 19728 21232 19780
rect 21548 19771 21600 19780
rect 21548 19737 21583 19771
rect 21583 19737 21600 19771
rect 21548 19728 21600 19737
rect 12808 19660 12860 19712
rect 14096 19660 14148 19712
rect 16120 19660 16172 19712
rect 16580 19660 16632 19712
rect 17776 19660 17828 19712
rect 20904 19703 20956 19712
rect 20904 19669 20913 19703
rect 20913 19669 20947 19703
rect 20947 19669 20956 19703
rect 20904 19660 20956 19669
rect 23296 19728 23348 19780
rect 4761 19558 4813 19610
rect 4825 19558 4877 19610
rect 4889 19558 4941 19610
rect 4953 19558 5005 19610
rect 5017 19558 5069 19610
rect 11063 19558 11115 19610
rect 11127 19558 11179 19610
rect 11191 19558 11243 19610
rect 11255 19558 11307 19610
rect 11319 19558 11371 19610
rect 17365 19558 17417 19610
rect 17429 19558 17481 19610
rect 17493 19558 17545 19610
rect 17557 19558 17609 19610
rect 17621 19558 17673 19610
rect 23667 19558 23719 19610
rect 23731 19558 23783 19610
rect 23795 19558 23847 19610
rect 23859 19558 23911 19610
rect 23923 19558 23975 19610
rect 2964 19456 3016 19508
rect 4436 19456 4488 19508
rect 1676 19431 1728 19440
rect 1676 19397 1685 19431
rect 1685 19397 1719 19431
rect 1719 19397 1728 19431
rect 1676 19388 1728 19397
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2780 19320 2832 19372
rect 4620 19388 4672 19440
rect 4804 19499 4856 19508
rect 4804 19465 4813 19499
rect 4813 19465 4847 19499
rect 4847 19465 4856 19499
rect 4804 19456 4856 19465
rect 8484 19456 8536 19508
rect 7196 19388 7248 19440
rect 9312 19388 9364 19440
rect 3148 19252 3200 19304
rect 5172 19320 5224 19372
rect 5816 19320 5868 19372
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 6736 19320 6788 19372
rect 8024 19320 8076 19372
rect 9496 19363 9548 19372
rect 9496 19329 9505 19363
rect 9505 19329 9539 19363
rect 9539 19329 9548 19363
rect 9496 19320 9548 19329
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 12716 19456 12768 19508
rect 14004 19499 14056 19508
rect 14004 19465 14013 19499
rect 14013 19465 14047 19499
rect 14047 19465 14056 19499
rect 14004 19456 14056 19465
rect 15200 19456 15252 19508
rect 12072 19388 12124 19440
rect 12808 19388 12860 19440
rect 13636 19431 13688 19440
rect 13636 19397 13645 19431
rect 13645 19397 13679 19431
rect 13679 19397 13688 19431
rect 13636 19388 13688 19397
rect 11520 19320 11572 19329
rect 3424 19159 3476 19168
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 3424 19116 3476 19125
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 4344 19252 4396 19304
rect 4436 19184 4488 19236
rect 12164 19252 12216 19304
rect 15752 19295 15804 19304
rect 15752 19261 15761 19295
rect 15761 19261 15795 19295
rect 15795 19261 15804 19295
rect 15752 19252 15804 19261
rect 15936 19320 15988 19372
rect 17132 19320 17184 19372
rect 17224 19252 17276 19304
rect 17868 19431 17920 19440
rect 17868 19397 17877 19431
rect 17877 19397 17911 19431
rect 17911 19397 17920 19431
rect 17868 19388 17920 19397
rect 17960 19388 18012 19440
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 18144 19320 18196 19372
rect 19156 19388 19208 19440
rect 19984 19388 20036 19440
rect 20168 19388 20220 19440
rect 20536 19456 20588 19508
rect 21272 19456 21324 19508
rect 23296 19456 23348 19508
rect 20720 19388 20772 19440
rect 20904 19388 20956 19440
rect 19340 19320 19392 19372
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 6000 19116 6052 19168
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 12624 19116 12676 19168
rect 14280 19116 14332 19168
rect 16580 19184 16632 19236
rect 17316 19227 17368 19236
rect 17316 19193 17325 19227
rect 17325 19193 17359 19227
rect 17359 19193 17368 19227
rect 17316 19184 17368 19193
rect 18512 19295 18564 19304
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 21088 19320 21140 19372
rect 21640 19388 21692 19440
rect 21824 19363 21876 19372
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 18144 19184 18196 19236
rect 18236 19184 18288 19236
rect 17040 19159 17092 19168
rect 17040 19125 17049 19159
rect 17049 19125 17083 19159
rect 17083 19125 17092 19159
rect 17040 19116 17092 19125
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17224 19116 17276 19125
rect 17408 19116 17460 19168
rect 20720 19295 20772 19304
rect 20720 19261 20729 19295
rect 20729 19261 20763 19295
rect 20763 19261 20772 19295
rect 20720 19252 20772 19261
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 23388 19320 23440 19372
rect 20444 19184 20496 19236
rect 21456 19184 21508 19236
rect 22008 19184 22060 19236
rect 21548 19116 21600 19168
rect 4101 19014 4153 19066
rect 4165 19014 4217 19066
rect 4229 19014 4281 19066
rect 4293 19014 4345 19066
rect 4357 19014 4409 19066
rect 10403 19014 10455 19066
rect 10467 19014 10519 19066
rect 10531 19014 10583 19066
rect 10595 19014 10647 19066
rect 10659 19014 10711 19066
rect 16705 19014 16757 19066
rect 16769 19014 16821 19066
rect 16833 19014 16885 19066
rect 16897 19014 16949 19066
rect 16961 19014 17013 19066
rect 23007 19014 23059 19066
rect 23071 19014 23123 19066
rect 23135 19014 23187 19066
rect 23199 19014 23251 19066
rect 23263 19014 23315 19066
rect 2780 18912 2832 18964
rect 6460 18912 6512 18964
rect 7196 18955 7248 18964
rect 7196 18921 7205 18955
rect 7205 18921 7239 18955
rect 7239 18921 7248 18955
rect 7196 18912 7248 18921
rect 9680 18912 9732 18964
rect 11428 18912 11480 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 14556 18912 14608 18964
rect 19248 18912 19300 18964
rect 19340 18912 19392 18964
rect 20076 18912 20128 18964
rect 20260 18955 20312 18964
rect 20260 18921 20269 18955
rect 20269 18921 20303 18955
rect 20303 18921 20312 18955
rect 20260 18912 20312 18921
rect 20628 18912 20680 18964
rect 20720 18912 20772 18964
rect 21088 18912 21140 18964
rect 14464 18887 14516 18896
rect 14464 18853 14473 18887
rect 14473 18853 14507 18887
rect 14507 18853 14516 18887
rect 14464 18844 14516 18853
rect 16488 18844 16540 18896
rect 17040 18844 17092 18896
rect 5264 18776 5316 18828
rect 5540 18776 5592 18828
rect 6368 18776 6420 18828
rect 10324 18819 10376 18828
rect 10324 18785 10333 18819
rect 10333 18785 10367 18819
rect 10367 18785 10376 18819
rect 10324 18776 10376 18785
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 6552 18708 6604 18760
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 11520 18708 11572 18760
rect 5264 18683 5316 18692
rect 5264 18649 5273 18683
rect 5273 18649 5307 18683
rect 5307 18649 5316 18683
rect 5264 18640 5316 18649
rect 11336 18640 11388 18692
rect 12992 18708 13044 18760
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 12716 18640 12768 18692
rect 14372 18708 14424 18760
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 16120 18708 16172 18760
rect 17316 18708 17368 18760
rect 17776 18708 17828 18760
rect 17960 18708 18012 18760
rect 20076 18819 20128 18828
rect 20076 18785 20085 18819
rect 20085 18785 20119 18819
rect 20119 18785 20128 18819
rect 20076 18776 20128 18785
rect 19616 18708 19668 18760
rect 13636 18640 13688 18692
rect 14188 18640 14240 18692
rect 14832 18640 14884 18692
rect 16396 18683 16448 18692
rect 16396 18649 16405 18683
rect 16405 18649 16439 18683
rect 16439 18649 16448 18683
rect 16396 18640 16448 18649
rect 5172 18572 5224 18624
rect 8760 18572 8812 18624
rect 10140 18615 10192 18624
rect 10140 18581 10149 18615
rect 10149 18581 10183 18615
rect 10183 18581 10192 18615
rect 10140 18572 10192 18581
rect 12900 18572 12952 18624
rect 15752 18572 15804 18624
rect 19800 18708 19852 18760
rect 20720 18708 20772 18760
rect 21088 18819 21140 18828
rect 21088 18785 21097 18819
rect 21097 18785 21131 18819
rect 21131 18785 21140 18819
rect 21088 18776 21140 18785
rect 23480 18844 23532 18896
rect 16856 18615 16908 18624
rect 16856 18581 16865 18615
rect 16865 18581 16899 18615
rect 16899 18581 16908 18615
rect 16856 18572 16908 18581
rect 17040 18572 17092 18624
rect 17224 18572 17276 18624
rect 17776 18615 17828 18624
rect 17776 18581 17785 18615
rect 17785 18581 17819 18615
rect 17819 18581 17828 18615
rect 17776 18572 17828 18581
rect 18236 18615 18288 18624
rect 18236 18581 18245 18615
rect 18245 18581 18279 18615
rect 18279 18581 18288 18615
rect 18236 18572 18288 18581
rect 18696 18615 18748 18624
rect 18696 18581 18705 18615
rect 18705 18581 18739 18615
rect 18739 18581 18748 18615
rect 18696 18572 18748 18581
rect 20536 18640 20588 18692
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 21364 18708 21416 18760
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 21456 18683 21508 18692
rect 21456 18649 21465 18683
rect 21465 18649 21499 18683
rect 21499 18649 21508 18683
rect 21456 18640 21508 18649
rect 21548 18683 21600 18692
rect 21548 18649 21557 18683
rect 21557 18649 21591 18683
rect 21591 18649 21600 18683
rect 21548 18640 21600 18649
rect 19800 18572 19852 18624
rect 20352 18572 20404 18624
rect 21088 18572 21140 18624
rect 4761 18470 4813 18522
rect 4825 18470 4877 18522
rect 4889 18470 4941 18522
rect 4953 18470 5005 18522
rect 5017 18470 5069 18522
rect 11063 18470 11115 18522
rect 11127 18470 11179 18522
rect 11191 18470 11243 18522
rect 11255 18470 11307 18522
rect 11319 18470 11371 18522
rect 17365 18470 17417 18522
rect 17429 18470 17481 18522
rect 17493 18470 17545 18522
rect 17557 18470 17609 18522
rect 17621 18470 17673 18522
rect 23667 18470 23719 18522
rect 23731 18470 23783 18522
rect 23795 18470 23847 18522
rect 23859 18470 23911 18522
rect 23923 18470 23975 18522
rect 3792 18368 3844 18420
rect 5264 18368 5316 18420
rect 8576 18411 8628 18420
rect 8576 18377 8585 18411
rect 8585 18377 8619 18411
rect 8619 18377 8628 18411
rect 8576 18368 8628 18377
rect 3240 18300 3292 18352
rect 9312 18300 9364 18352
rect 3056 18207 3108 18216
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 3056 18164 3108 18173
rect 3608 18164 3660 18216
rect 4436 18207 4488 18216
rect 4436 18173 4445 18207
rect 4445 18173 4479 18207
rect 4479 18173 4488 18207
rect 4436 18164 4488 18173
rect 4712 18275 4764 18284
rect 4712 18241 4721 18275
rect 4721 18241 4755 18275
rect 4755 18241 4764 18275
rect 4712 18232 4764 18241
rect 5080 18164 5132 18216
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 4528 18096 4580 18148
rect 5448 18207 5500 18216
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 6000 18275 6052 18284
rect 6000 18241 6009 18275
rect 6009 18241 6043 18275
rect 6043 18241 6052 18275
rect 6000 18232 6052 18241
rect 6184 18275 6236 18284
rect 6184 18241 6193 18275
rect 6193 18241 6227 18275
rect 6227 18241 6236 18275
rect 6184 18232 6236 18241
rect 10784 18368 10836 18420
rect 11888 18368 11940 18420
rect 10324 18300 10376 18352
rect 6828 18164 6880 18216
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 5632 18096 5684 18148
rect 9956 18164 10008 18216
rect 10784 18275 10836 18284
rect 10784 18241 10793 18275
rect 10793 18241 10827 18275
rect 10827 18241 10836 18275
rect 10784 18232 10836 18241
rect 10876 18275 10928 18284
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 11060 18275 11112 18284
rect 11060 18241 11069 18275
rect 11069 18241 11103 18275
rect 11103 18241 11112 18275
rect 11060 18232 11112 18241
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 11888 18275 11940 18284
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 12624 18232 12676 18284
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 13912 18275 13964 18284
rect 13912 18241 13921 18275
rect 13921 18241 13955 18275
rect 13955 18241 13964 18275
rect 13912 18232 13964 18241
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 14556 18368 14608 18420
rect 15936 18368 15988 18420
rect 16948 18368 17000 18420
rect 17960 18411 18012 18420
rect 17960 18377 17995 18411
rect 17995 18377 18012 18411
rect 17960 18368 18012 18377
rect 18696 18368 18748 18420
rect 19708 18368 19760 18420
rect 20168 18411 20220 18420
rect 20168 18377 20177 18411
rect 20177 18377 20211 18411
rect 20211 18377 20220 18411
rect 20168 18368 20220 18377
rect 16120 18343 16172 18352
rect 16120 18309 16129 18343
rect 16129 18309 16163 18343
rect 16163 18309 16172 18343
rect 16120 18300 16172 18309
rect 14648 18275 14700 18284
rect 14648 18241 14657 18275
rect 14657 18241 14691 18275
rect 14691 18241 14700 18275
rect 14648 18232 14700 18241
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 18144 18300 18196 18352
rect 19800 18343 19852 18352
rect 19800 18309 19809 18343
rect 19809 18309 19843 18343
rect 19843 18309 19852 18343
rect 19800 18300 19852 18309
rect 20352 18300 20404 18352
rect 21364 18411 21416 18420
rect 21364 18377 21373 18411
rect 21373 18377 21407 18411
rect 21407 18377 21416 18411
rect 21364 18368 21416 18377
rect 25136 18411 25188 18420
rect 25136 18377 25145 18411
rect 25145 18377 25179 18411
rect 25179 18377 25188 18411
rect 25136 18368 25188 18377
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 18236 18232 18288 18284
rect 20720 18232 20772 18284
rect 20996 18275 21048 18284
rect 20996 18241 21005 18275
rect 21005 18241 21039 18275
rect 21039 18241 21048 18275
rect 20996 18232 21048 18241
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 21456 18300 21508 18352
rect 1676 18028 1728 18080
rect 3608 18071 3660 18080
rect 3608 18037 3617 18071
rect 3617 18037 3651 18071
rect 3651 18037 3660 18071
rect 3608 18028 3660 18037
rect 4804 18071 4856 18080
rect 4804 18037 4813 18071
rect 4813 18037 4847 18071
rect 4847 18037 4856 18071
rect 4804 18028 4856 18037
rect 5356 18071 5408 18080
rect 5356 18037 5365 18071
rect 5365 18037 5399 18071
rect 5399 18037 5408 18071
rect 5356 18028 5408 18037
rect 5448 18028 5500 18080
rect 9036 18071 9088 18080
rect 9036 18037 9045 18071
rect 9045 18037 9079 18071
rect 9079 18037 9088 18071
rect 9036 18028 9088 18037
rect 10784 18028 10836 18080
rect 11336 18028 11388 18080
rect 11704 18028 11756 18080
rect 13084 18096 13136 18148
rect 12992 18028 13044 18080
rect 16488 18139 16540 18148
rect 16488 18105 16497 18139
rect 16497 18105 16531 18139
rect 16531 18105 16540 18139
rect 20628 18164 20680 18216
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 16488 18096 16540 18105
rect 17224 18096 17276 18148
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 14556 18071 14608 18080
rect 14556 18037 14565 18071
rect 14565 18037 14599 18071
rect 14599 18037 14608 18071
rect 14556 18028 14608 18037
rect 15016 18028 15068 18080
rect 16212 18028 16264 18080
rect 16948 18028 17000 18080
rect 20444 18096 20496 18148
rect 20996 18096 21048 18148
rect 17408 18028 17460 18080
rect 19800 18028 19852 18080
rect 20260 18028 20312 18080
rect 4101 17926 4153 17978
rect 4165 17926 4217 17978
rect 4229 17926 4281 17978
rect 4293 17926 4345 17978
rect 4357 17926 4409 17978
rect 10403 17926 10455 17978
rect 10467 17926 10519 17978
rect 10531 17926 10583 17978
rect 10595 17926 10647 17978
rect 10659 17926 10711 17978
rect 16705 17926 16757 17978
rect 16769 17926 16821 17978
rect 16833 17926 16885 17978
rect 16897 17926 16949 17978
rect 16961 17926 17013 17978
rect 23007 17926 23059 17978
rect 23071 17926 23123 17978
rect 23135 17926 23187 17978
rect 23199 17926 23251 17978
rect 23263 17926 23315 17978
rect 4804 17824 4856 17876
rect 5724 17824 5776 17876
rect 6460 17824 6512 17876
rect 6736 17824 6788 17876
rect 7472 17824 7524 17876
rect 6184 17756 6236 17808
rect 7380 17799 7432 17808
rect 7380 17765 7389 17799
rect 7389 17765 7423 17799
rect 7423 17765 7432 17799
rect 7380 17756 7432 17765
rect 8392 17756 8444 17808
rect 10232 17756 10284 17808
rect 10876 17756 10928 17808
rect 11888 17756 11940 17808
rect 4436 17688 4488 17740
rect 5080 17688 5132 17740
rect 5540 17688 5592 17740
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 3056 17620 3108 17672
rect 3332 17620 3384 17672
rect 5172 17620 5224 17672
rect 5356 17620 5408 17672
rect 1676 17595 1728 17604
rect 1676 17561 1685 17595
rect 1685 17561 1719 17595
rect 1719 17561 1728 17595
rect 1676 17552 1728 17561
rect 2412 17552 2464 17604
rect 3608 17552 3660 17604
rect 4712 17484 4764 17536
rect 12072 17731 12124 17740
rect 12072 17697 12081 17731
rect 12081 17697 12115 17731
rect 12115 17697 12124 17731
rect 12072 17688 12124 17697
rect 13176 17824 13228 17876
rect 13912 17824 13964 17876
rect 14280 17867 14332 17876
rect 14280 17833 14289 17867
rect 14289 17833 14323 17867
rect 14323 17833 14332 17867
rect 14280 17824 14332 17833
rect 17040 17824 17092 17876
rect 13820 17756 13872 17808
rect 16120 17688 16172 17740
rect 6000 17620 6052 17672
rect 6644 17620 6696 17672
rect 6828 17663 6880 17672
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 7104 17663 7156 17672
rect 7104 17629 7113 17663
rect 7113 17629 7147 17663
rect 7147 17629 7156 17663
rect 7104 17620 7156 17629
rect 9128 17620 9180 17672
rect 7288 17552 7340 17604
rect 10140 17595 10192 17604
rect 10140 17561 10149 17595
rect 10149 17561 10183 17595
rect 10183 17561 10192 17595
rect 10140 17552 10192 17561
rect 12440 17620 12492 17672
rect 13728 17620 13780 17672
rect 18144 17756 18196 17808
rect 11520 17552 11572 17604
rect 11796 17552 11848 17604
rect 12900 17595 12952 17604
rect 12900 17561 12909 17595
rect 12909 17561 12943 17595
rect 12943 17561 12952 17595
rect 12900 17552 12952 17561
rect 13360 17595 13412 17604
rect 13360 17561 13369 17595
rect 13369 17561 13403 17595
rect 13403 17561 13412 17595
rect 13360 17552 13412 17561
rect 13544 17595 13596 17604
rect 13544 17561 13553 17595
rect 13553 17561 13587 17595
rect 13587 17561 13596 17595
rect 13544 17552 13596 17561
rect 14188 17552 14240 17604
rect 5632 17484 5684 17536
rect 6000 17484 6052 17536
rect 6184 17484 6236 17536
rect 6276 17527 6328 17536
rect 6276 17493 6285 17527
rect 6285 17493 6319 17527
rect 6319 17493 6328 17527
rect 6276 17484 6328 17493
rect 6644 17484 6696 17536
rect 7932 17527 7984 17536
rect 7932 17493 7941 17527
rect 7941 17493 7975 17527
rect 7975 17493 7984 17527
rect 7932 17484 7984 17493
rect 8668 17484 8720 17536
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 8760 17484 8812 17493
rect 8944 17484 8996 17536
rect 11428 17484 11480 17536
rect 12532 17484 12584 17536
rect 13912 17484 13964 17536
rect 17132 17620 17184 17672
rect 17960 17688 18012 17740
rect 20076 17688 20128 17740
rect 20260 17688 20312 17740
rect 23480 17731 23532 17740
rect 14740 17527 14792 17536
rect 14740 17493 14749 17527
rect 14749 17493 14783 17527
rect 14783 17493 14792 17527
rect 14740 17484 14792 17493
rect 14832 17484 14884 17536
rect 18236 17552 18288 17604
rect 19616 17620 19668 17672
rect 19892 17620 19944 17672
rect 20536 17620 20588 17672
rect 21180 17620 21232 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 23480 17697 23489 17731
rect 23489 17697 23523 17731
rect 23523 17697 23532 17731
rect 23480 17688 23532 17697
rect 23388 17620 23440 17672
rect 19984 17552 20036 17604
rect 20720 17552 20772 17604
rect 21364 17595 21416 17604
rect 21364 17561 21373 17595
rect 21373 17561 21407 17595
rect 21407 17561 21416 17595
rect 21364 17552 21416 17561
rect 18420 17484 18472 17536
rect 19708 17484 19760 17536
rect 20076 17484 20128 17536
rect 22284 17484 22336 17536
rect 22744 17527 22796 17536
rect 22744 17493 22753 17527
rect 22753 17493 22787 17527
rect 22787 17493 22796 17527
rect 22744 17484 22796 17493
rect 4761 17382 4813 17434
rect 4825 17382 4877 17434
rect 4889 17382 4941 17434
rect 4953 17382 5005 17434
rect 5017 17382 5069 17434
rect 11063 17382 11115 17434
rect 11127 17382 11179 17434
rect 11191 17382 11243 17434
rect 11255 17382 11307 17434
rect 11319 17382 11371 17434
rect 17365 17382 17417 17434
rect 17429 17382 17481 17434
rect 17493 17382 17545 17434
rect 17557 17382 17609 17434
rect 17621 17382 17673 17434
rect 23667 17382 23719 17434
rect 23731 17382 23783 17434
rect 23795 17382 23847 17434
rect 23859 17382 23911 17434
rect 23923 17382 23975 17434
rect 2412 17280 2464 17332
rect 7472 17280 7524 17332
rect 6184 17212 6236 17264
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 2320 17144 2372 17196
rect 4436 17187 4488 17196
rect 4436 17153 4445 17187
rect 4445 17153 4479 17187
rect 4479 17153 4488 17187
rect 4436 17144 4488 17153
rect 6000 17144 6052 17196
rect 6460 17212 6512 17264
rect 9312 17323 9364 17332
rect 9312 17289 9321 17323
rect 9321 17289 9355 17323
rect 9355 17289 9364 17323
rect 9312 17280 9364 17289
rect 10140 17280 10192 17332
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 5724 17008 5776 17060
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 6552 17076 6604 17128
rect 8944 17144 8996 17196
rect 9772 17212 9824 17264
rect 7012 17076 7064 17128
rect 9036 17076 9088 17128
rect 9312 17076 9364 17128
rect 10324 17144 10376 17196
rect 9956 17008 10008 17060
rect 5356 16940 5408 16992
rect 6368 16940 6420 16992
rect 6736 16983 6788 16992
rect 6736 16949 6745 16983
rect 6745 16949 6779 16983
rect 6779 16949 6788 16983
rect 6736 16940 6788 16949
rect 6828 16940 6880 16992
rect 8944 16940 8996 16992
rect 10232 16940 10284 16992
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 11612 17144 11664 17196
rect 14740 17280 14792 17332
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 11888 17119 11940 17128
rect 11888 17085 11897 17119
rect 11897 17085 11931 17119
rect 11931 17085 11940 17119
rect 11888 17076 11940 17085
rect 12716 17076 12768 17128
rect 14004 17212 14056 17264
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 18236 17280 18288 17332
rect 18420 17323 18472 17332
rect 18420 17289 18429 17323
rect 18429 17289 18463 17323
rect 18463 17289 18472 17323
rect 18420 17280 18472 17289
rect 21272 17280 21324 17332
rect 17960 17212 18012 17264
rect 14188 17076 14240 17128
rect 19800 17144 19852 17196
rect 22284 17255 22336 17264
rect 22284 17221 22293 17255
rect 22293 17221 22327 17255
rect 22327 17221 22336 17255
rect 22284 17212 22336 17221
rect 13636 17008 13688 17060
rect 16580 17076 16632 17128
rect 19984 17119 20036 17128
rect 19984 17085 19993 17119
rect 19993 17085 20027 17119
rect 20027 17085 20036 17119
rect 19984 17076 20036 17085
rect 20536 17119 20588 17128
rect 20536 17085 20545 17119
rect 20545 17085 20579 17119
rect 20579 17085 20588 17119
rect 20536 17076 20588 17085
rect 21456 17144 21508 17196
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 25688 17187 25740 17196
rect 25688 17153 25697 17187
rect 25697 17153 25731 17187
rect 25731 17153 25740 17187
rect 25688 17144 25740 17153
rect 20996 17119 21048 17128
rect 20996 17085 21005 17119
rect 21005 17085 21039 17119
rect 21039 17085 21048 17119
rect 20996 17076 21048 17085
rect 23480 17076 23532 17128
rect 20076 17008 20128 17060
rect 25872 17051 25924 17060
rect 25872 17017 25881 17051
rect 25881 17017 25915 17051
rect 25915 17017 25924 17051
rect 25872 17008 25924 17017
rect 10876 16940 10928 16992
rect 14188 16940 14240 16992
rect 14648 16940 14700 16992
rect 15108 16940 15160 16992
rect 18512 16940 18564 16992
rect 20904 16940 20956 16992
rect 4101 16838 4153 16890
rect 4165 16838 4217 16890
rect 4229 16838 4281 16890
rect 4293 16838 4345 16890
rect 4357 16838 4409 16890
rect 10403 16838 10455 16890
rect 10467 16838 10519 16890
rect 10531 16838 10583 16890
rect 10595 16838 10647 16890
rect 10659 16838 10711 16890
rect 16705 16838 16757 16890
rect 16769 16838 16821 16890
rect 16833 16838 16885 16890
rect 16897 16838 16949 16890
rect 16961 16838 17013 16890
rect 23007 16838 23059 16890
rect 23071 16838 23123 16890
rect 23135 16838 23187 16890
rect 23199 16838 23251 16890
rect 23263 16838 23315 16890
rect 2136 16736 2188 16788
rect 4620 16779 4672 16788
rect 4620 16745 4629 16779
rect 4629 16745 4663 16779
rect 4663 16745 4672 16779
rect 4620 16736 4672 16745
rect 4712 16736 4764 16788
rect 6092 16736 6144 16788
rect 6828 16736 6880 16788
rect 940 16532 992 16584
rect 6460 16668 6512 16720
rect 5816 16600 5868 16652
rect 6276 16600 6328 16652
rect 6552 16600 6604 16652
rect 8668 16736 8720 16788
rect 9128 16668 9180 16720
rect 9956 16668 10008 16720
rect 10048 16668 10100 16720
rect 3976 16396 4028 16448
rect 5724 16532 5776 16584
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 10324 16600 10376 16652
rect 9128 16532 9180 16584
rect 9772 16575 9824 16584
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 7288 16507 7340 16516
rect 7288 16473 7297 16507
rect 7297 16473 7331 16507
rect 7331 16473 7340 16507
rect 7288 16464 7340 16473
rect 5540 16396 5592 16448
rect 6644 16396 6696 16448
rect 10324 16507 10376 16516
rect 10324 16473 10333 16507
rect 10333 16473 10367 16507
rect 10367 16473 10376 16507
rect 10324 16464 10376 16473
rect 11336 16600 11388 16652
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 12072 16668 12124 16720
rect 14004 16736 14056 16788
rect 13636 16668 13688 16720
rect 18512 16668 18564 16720
rect 13452 16600 13504 16652
rect 14372 16600 14424 16652
rect 20720 16736 20772 16788
rect 20904 16736 20956 16788
rect 25688 16736 25740 16788
rect 20812 16668 20864 16720
rect 23204 16711 23256 16720
rect 23204 16677 23213 16711
rect 23213 16677 23247 16711
rect 23247 16677 23256 16711
rect 23204 16668 23256 16677
rect 15568 16532 15620 16584
rect 12440 16507 12492 16516
rect 12440 16473 12449 16507
rect 12449 16473 12483 16507
rect 12483 16473 12492 16507
rect 12440 16464 12492 16473
rect 17960 16532 18012 16584
rect 19892 16600 19944 16652
rect 18052 16464 18104 16516
rect 12072 16396 12124 16448
rect 20260 16575 20312 16584
rect 20260 16541 20269 16575
rect 20269 16541 20303 16575
rect 20303 16541 20312 16575
rect 20260 16532 20312 16541
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20536 16532 20588 16541
rect 20720 16575 20772 16584
rect 20720 16541 20729 16575
rect 20729 16541 20763 16575
rect 20763 16541 20772 16575
rect 20720 16532 20772 16541
rect 21364 16600 21416 16652
rect 21456 16643 21508 16652
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 22100 16600 22152 16652
rect 20168 16464 20220 16516
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 23572 16600 23624 16652
rect 20996 16507 21048 16516
rect 20996 16473 21005 16507
rect 21005 16473 21039 16507
rect 21039 16473 21048 16507
rect 20996 16464 21048 16473
rect 21824 16464 21876 16516
rect 22744 16464 22796 16516
rect 21088 16439 21140 16448
rect 21088 16405 21103 16439
rect 21103 16405 21137 16439
rect 21137 16405 21140 16439
rect 21088 16396 21140 16405
rect 23480 16439 23532 16448
rect 23480 16405 23489 16439
rect 23489 16405 23523 16439
rect 23523 16405 23532 16439
rect 23480 16396 23532 16405
rect 4761 16294 4813 16346
rect 4825 16294 4877 16346
rect 4889 16294 4941 16346
rect 4953 16294 5005 16346
rect 5017 16294 5069 16346
rect 11063 16294 11115 16346
rect 11127 16294 11179 16346
rect 11191 16294 11243 16346
rect 11255 16294 11307 16346
rect 11319 16294 11371 16346
rect 17365 16294 17417 16346
rect 17429 16294 17481 16346
rect 17493 16294 17545 16346
rect 17557 16294 17609 16346
rect 17621 16294 17673 16346
rect 23667 16294 23719 16346
rect 23731 16294 23783 16346
rect 23795 16294 23847 16346
rect 23859 16294 23911 16346
rect 23923 16294 23975 16346
rect 2320 16192 2372 16244
rect 3792 16192 3844 16244
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 5448 16124 5500 16176
rect 6644 16192 6696 16244
rect 7288 16192 7340 16244
rect 10324 16192 10376 16244
rect 11520 16192 11572 16244
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 13452 16235 13504 16244
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 8576 16124 8628 16176
rect 15108 16124 15160 16176
rect 3884 15988 3936 16040
rect 3976 16031 4028 16040
rect 3976 15997 3985 16031
rect 3985 15997 4019 16031
rect 4019 15997 4028 16031
rect 3976 15988 4028 15997
rect 2780 15920 2832 15972
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 9772 16056 9824 16108
rect 10784 16056 10836 16108
rect 1676 15852 1728 15904
rect 2228 15852 2280 15904
rect 2964 15852 3016 15904
rect 5172 15852 5224 15904
rect 6736 15920 6788 15972
rect 7564 16031 7616 16040
rect 7564 15997 7573 16031
rect 7573 15997 7607 16031
rect 7607 15997 7616 16031
rect 7564 15988 7616 15997
rect 10876 15988 10928 16040
rect 12532 16099 12584 16108
rect 12532 16065 12541 16099
rect 12541 16065 12575 16099
rect 12575 16065 12584 16099
rect 12532 16056 12584 16065
rect 16580 16056 16632 16108
rect 19248 16192 19300 16244
rect 20720 16192 20772 16244
rect 21180 16192 21232 16244
rect 18236 16124 18288 16176
rect 19064 16167 19116 16176
rect 19064 16133 19073 16167
rect 19073 16133 19107 16167
rect 19107 16133 19116 16167
rect 19064 16124 19116 16133
rect 21088 16124 21140 16176
rect 20812 16056 20864 16108
rect 12716 15988 12768 16040
rect 14648 15988 14700 16040
rect 17776 15988 17828 16040
rect 6000 15852 6052 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 17040 15852 17092 15904
rect 20996 16031 21048 16040
rect 20996 15997 21005 16031
rect 21005 15997 21039 16031
rect 21039 15997 21048 16031
rect 20996 15988 21048 15997
rect 21272 15988 21324 16040
rect 21824 15963 21876 15972
rect 21824 15929 21833 15963
rect 21833 15929 21867 15963
rect 21867 15929 21876 15963
rect 21824 15920 21876 15929
rect 4101 15750 4153 15802
rect 4165 15750 4217 15802
rect 4229 15750 4281 15802
rect 4293 15750 4345 15802
rect 4357 15750 4409 15802
rect 10403 15750 10455 15802
rect 10467 15750 10519 15802
rect 10531 15750 10583 15802
rect 10595 15750 10647 15802
rect 10659 15750 10711 15802
rect 16705 15750 16757 15802
rect 16769 15750 16821 15802
rect 16833 15750 16885 15802
rect 16897 15750 16949 15802
rect 16961 15750 17013 15802
rect 23007 15750 23059 15802
rect 23071 15750 23123 15802
rect 23135 15750 23187 15802
rect 23199 15750 23251 15802
rect 23263 15750 23315 15802
rect 2320 15648 2372 15700
rect 6000 15648 6052 15700
rect 7932 15648 7984 15700
rect 12440 15648 12492 15700
rect 17592 15648 17644 15700
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 18236 15648 18288 15700
rect 20996 15648 21048 15700
rect 3884 15580 3936 15632
rect 6460 15580 6512 15632
rect 13728 15580 13780 15632
rect 19064 15580 19116 15632
rect 1400 15512 1452 15564
rect 2228 15512 2280 15564
rect 4528 15512 4580 15564
rect 7380 15512 7432 15564
rect 2964 15444 3016 15496
rect 3792 15444 3844 15496
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 15476 15512 15528 15564
rect 15936 15512 15988 15564
rect 16948 15512 17000 15564
rect 17040 15512 17092 15564
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 7932 15487 7984 15496
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 7932 15444 7984 15453
rect 8116 15444 8168 15496
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 9956 15444 10008 15496
rect 11888 15444 11940 15496
rect 14464 15444 14516 15496
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 16488 15444 16540 15496
rect 19984 15512 20036 15564
rect 20628 15512 20680 15564
rect 21456 15512 21508 15564
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 19156 15444 19208 15496
rect 8576 15376 8628 15428
rect 17040 15376 17092 15428
rect 17868 15376 17920 15428
rect 4528 15308 4580 15360
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 7288 15308 7340 15360
rect 8300 15308 8352 15360
rect 9312 15308 9364 15360
rect 9772 15308 9824 15360
rect 10140 15351 10192 15360
rect 10140 15317 10149 15351
rect 10149 15317 10183 15351
rect 10183 15317 10192 15351
rect 10140 15308 10192 15317
rect 10232 15308 10284 15360
rect 13636 15308 13688 15360
rect 15752 15308 15804 15360
rect 16856 15308 16908 15360
rect 17684 15308 17736 15360
rect 20812 15444 20864 15496
rect 21088 15376 21140 15428
rect 23388 15308 23440 15360
rect 24308 15308 24360 15360
rect 4761 15206 4813 15258
rect 4825 15206 4877 15258
rect 4889 15206 4941 15258
rect 4953 15206 5005 15258
rect 5017 15206 5069 15258
rect 11063 15206 11115 15258
rect 11127 15206 11179 15258
rect 11191 15206 11243 15258
rect 11255 15206 11307 15258
rect 11319 15206 11371 15258
rect 17365 15206 17417 15258
rect 17429 15206 17481 15258
rect 17493 15206 17545 15258
rect 17557 15206 17609 15258
rect 17621 15206 17673 15258
rect 23667 15206 23719 15258
rect 23731 15206 23783 15258
rect 23795 15206 23847 15258
rect 23859 15206 23911 15258
rect 23923 15206 23975 15258
rect 1400 15104 1452 15156
rect 1676 15079 1728 15088
rect 1676 15045 1685 15079
rect 1685 15045 1719 15079
rect 1719 15045 1728 15079
rect 1676 15036 1728 15045
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 2780 14968 2832 15020
rect 5724 15036 5776 15088
rect 6552 15104 6604 15156
rect 7564 15104 7616 15156
rect 8116 15147 8168 15156
rect 8116 15113 8125 15147
rect 8125 15113 8159 15147
rect 8159 15113 8168 15147
rect 8116 15104 8168 15113
rect 7104 15036 7156 15088
rect 4896 14900 4948 14952
rect 5448 14900 5500 14952
rect 6644 14943 6696 14952
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 6644 14900 6696 14909
rect 6736 14900 6788 14952
rect 8576 15036 8628 15088
rect 9772 15036 9824 15088
rect 10140 15036 10192 15088
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 12164 15104 12216 15156
rect 12624 15079 12676 15088
rect 12624 15045 12633 15079
rect 12633 15045 12667 15079
rect 12667 15045 12676 15079
rect 12624 15036 12676 15045
rect 13728 15104 13780 15156
rect 16856 15104 16908 15156
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 21088 15104 21140 15156
rect 15752 15036 15804 15088
rect 17132 15036 17184 15088
rect 10784 14968 10836 15020
rect 8852 14943 8904 14952
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 7656 14832 7708 14884
rect 4528 14764 4580 14816
rect 9864 14764 9916 14816
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 11336 14900 11388 14952
rect 11796 14900 11848 14952
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 17316 14968 17368 15020
rect 12072 14900 12124 14952
rect 14740 14943 14792 14952
rect 14740 14909 14749 14943
rect 14749 14909 14783 14943
rect 14783 14909 14792 14943
rect 14740 14900 14792 14909
rect 18052 15011 18104 15020
rect 18052 14977 18061 15011
rect 18061 14977 18095 15011
rect 18095 14977 18104 15011
rect 18052 14968 18104 14977
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 18144 14900 18196 14952
rect 12624 14832 12676 14884
rect 18328 14832 18380 14884
rect 12256 14764 12308 14816
rect 12440 14764 12492 14816
rect 17960 14764 18012 14816
rect 18512 14764 18564 14816
rect 20076 14807 20128 14816
rect 20076 14773 20085 14807
rect 20085 14773 20119 14807
rect 20119 14773 20128 14807
rect 20076 14764 20128 14773
rect 20260 14764 20312 14816
rect 4101 14662 4153 14714
rect 4165 14662 4217 14714
rect 4229 14662 4281 14714
rect 4293 14662 4345 14714
rect 4357 14662 4409 14714
rect 10403 14662 10455 14714
rect 10467 14662 10519 14714
rect 10531 14662 10583 14714
rect 10595 14662 10647 14714
rect 10659 14662 10711 14714
rect 16705 14662 16757 14714
rect 16769 14662 16821 14714
rect 16833 14662 16885 14714
rect 16897 14662 16949 14714
rect 16961 14662 17013 14714
rect 23007 14662 23059 14714
rect 23071 14662 23123 14714
rect 23135 14662 23187 14714
rect 23199 14662 23251 14714
rect 23263 14662 23315 14714
rect 4896 14603 4948 14612
rect 4896 14569 4905 14603
rect 4905 14569 4939 14603
rect 4939 14569 4948 14603
rect 4896 14560 4948 14569
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 6644 14560 6696 14612
rect 7104 14560 7156 14612
rect 12532 14560 12584 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 14464 14603 14516 14612
rect 14464 14569 14473 14603
rect 14473 14569 14507 14603
rect 14507 14569 14516 14603
rect 14464 14560 14516 14569
rect 16304 14560 16356 14612
rect 17224 14603 17276 14612
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 6552 14492 6604 14544
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 11888 14492 11940 14544
rect 10876 14424 10928 14476
rect 11612 14424 11664 14476
rect 12072 14424 12124 14476
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 12808 14424 12860 14476
rect 15200 14492 15252 14544
rect 4528 14356 4580 14408
rect 5172 14356 5224 14408
rect 6000 14356 6052 14408
rect 6368 14356 6420 14408
rect 6828 14356 6880 14408
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 1952 14288 2004 14340
rect 5540 14288 5592 14340
rect 4620 14220 4672 14272
rect 5908 14220 5960 14272
rect 6736 14220 6788 14272
rect 7380 14288 7432 14340
rect 8300 14288 8352 14340
rect 8668 14220 8720 14272
rect 10232 14288 10284 14340
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 16580 14492 16632 14544
rect 18144 14560 18196 14612
rect 14372 14356 14424 14408
rect 17132 14356 17184 14408
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17868 14492 17920 14544
rect 12348 14288 12400 14340
rect 11520 14220 11572 14272
rect 13452 14220 13504 14272
rect 14280 14331 14332 14340
rect 14280 14297 14289 14331
rect 14289 14297 14323 14331
rect 14323 14297 14332 14331
rect 14280 14288 14332 14297
rect 14740 14288 14792 14340
rect 15200 14263 15252 14272
rect 15752 14331 15804 14340
rect 15752 14297 15761 14331
rect 15761 14297 15795 14331
rect 15795 14297 15804 14331
rect 15752 14288 15804 14297
rect 15936 14331 15988 14340
rect 15936 14297 15945 14331
rect 15945 14297 15979 14331
rect 15979 14297 15988 14331
rect 15936 14288 15988 14297
rect 16212 14331 16264 14340
rect 16212 14297 16221 14331
rect 16221 14297 16255 14331
rect 16255 14297 16264 14331
rect 16212 14288 16264 14297
rect 15200 14229 15215 14263
rect 15215 14229 15249 14263
rect 15249 14229 15252 14263
rect 15200 14220 15252 14229
rect 18144 14356 18196 14408
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 19248 14467 19300 14476
rect 19248 14433 19257 14467
rect 19257 14433 19291 14467
rect 19291 14433 19300 14467
rect 19248 14424 19300 14433
rect 18972 14399 19024 14408
rect 18972 14365 18981 14399
rect 18981 14365 19015 14399
rect 19015 14365 19024 14399
rect 18972 14356 19024 14365
rect 19432 14288 19484 14340
rect 20076 14288 20128 14340
rect 20168 14220 20220 14272
rect 4761 14118 4813 14170
rect 4825 14118 4877 14170
rect 4889 14118 4941 14170
rect 4953 14118 5005 14170
rect 5017 14118 5069 14170
rect 11063 14118 11115 14170
rect 11127 14118 11179 14170
rect 11191 14118 11243 14170
rect 11255 14118 11307 14170
rect 11319 14118 11371 14170
rect 17365 14118 17417 14170
rect 17429 14118 17481 14170
rect 17493 14118 17545 14170
rect 17557 14118 17609 14170
rect 17621 14118 17673 14170
rect 23667 14118 23719 14170
rect 23731 14118 23783 14170
rect 23795 14118 23847 14170
rect 23859 14118 23911 14170
rect 23923 14118 23975 14170
rect 4620 13948 4672 14000
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 6828 14016 6880 14068
rect 7380 14059 7432 14068
rect 7380 14025 7389 14059
rect 7389 14025 7423 14059
rect 7423 14025 7432 14059
rect 7380 14016 7432 14025
rect 9128 14016 9180 14068
rect 9496 14016 9548 14068
rect 3884 13812 3936 13864
rect 5908 13923 5960 13932
rect 5908 13889 5917 13923
rect 5917 13889 5951 13923
rect 5951 13889 5960 13923
rect 5908 13880 5960 13889
rect 7472 13948 7524 14000
rect 7656 13948 7708 14000
rect 8668 13948 8720 14000
rect 10048 13948 10100 14000
rect 10784 13948 10836 14000
rect 11520 14016 11572 14068
rect 11796 14016 11848 14068
rect 11980 14016 12032 14068
rect 12256 14016 12308 14068
rect 12808 14016 12860 14068
rect 12900 14016 12952 14068
rect 17132 14016 17184 14068
rect 17500 14016 17552 14068
rect 18972 14016 19024 14068
rect 11888 13948 11940 14000
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 7196 13880 7248 13932
rect 7288 13880 7340 13932
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 10324 13880 10376 13932
rect 13636 13880 13688 13932
rect 14372 13880 14424 13932
rect 6736 13744 6788 13796
rect 8760 13744 8812 13796
rect 9496 13812 9548 13864
rect 10876 13812 10928 13864
rect 11704 13744 11756 13796
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 14464 13812 14516 13864
rect 15752 13812 15804 13864
rect 16304 13812 16356 13864
rect 16948 13812 17000 13864
rect 17224 13991 17276 14000
rect 17224 13957 17249 13991
rect 17249 13957 17276 13991
rect 17224 13948 17276 13957
rect 17592 13991 17644 14000
rect 17592 13957 17601 13991
rect 17601 13957 17635 13991
rect 17635 13957 17644 13991
rect 17592 13948 17644 13957
rect 17224 13812 17276 13864
rect 18052 13948 18104 14000
rect 18696 13948 18748 14000
rect 20260 13948 20312 14000
rect 19156 13880 19208 13932
rect 17868 13744 17920 13796
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 5908 13676 5960 13728
rect 6092 13719 6144 13728
rect 6092 13685 6101 13719
rect 6101 13685 6135 13719
rect 6135 13685 6144 13719
rect 6092 13676 6144 13685
rect 7380 13676 7432 13728
rect 11520 13676 11572 13728
rect 11796 13676 11848 13728
rect 16488 13676 16540 13728
rect 19800 13812 19852 13864
rect 18880 13744 18932 13796
rect 20352 13676 20404 13728
rect 4101 13574 4153 13626
rect 4165 13574 4217 13626
rect 4229 13574 4281 13626
rect 4293 13574 4345 13626
rect 4357 13574 4409 13626
rect 10403 13574 10455 13626
rect 10467 13574 10519 13626
rect 10531 13574 10583 13626
rect 10595 13574 10647 13626
rect 10659 13574 10711 13626
rect 16705 13574 16757 13626
rect 16769 13574 16821 13626
rect 16833 13574 16885 13626
rect 16897 13574 16949 13626
rect 16961 13574 17013 13626
rect 23007 13574 23059 13626
rect 23071 13574 23123 13626
rect 23135 13574 23187 13626
rect 23199 13574 23251 13626
rect 23263 13574 23315 13626
rect 5908 13472 5960 13524
rect 6736 13515 6788 13524
rect 6736 13481 6745 13515
rect 6745 13481 6779 13515
rect 6779 13481 6788 13515
rect 6736 13472 6788 13481
rect 7012 13472 7064 13524
rect 12624 13472 12676 13524
rect 15936 13472 15988 13524
rect 17776 13472 17828 13524
rect 17960 13472 18012 13524
rect 5264 13404 5316 13456
rect 6092 13336 6144 13388
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 5172 13268 5224 13320
rect 6184 13268 6236 13320
rect 7196 13336 7248 13388
rect 16304 13447 16356 13456
rect 16304 13413 16313 13447
rect 16313 13413 16347 13447
rect 16347 13413 16356 13447
rect 16304 13404 16356 13413
rect 11612 13336 11664 13388
rect 7656 13268 7708 13320
rect 10876 13268 10928 13320
rect 13452 13336 13504 13388
rect 11796 13268 11848 13320
rect 12348 13311 12400 13320
rect 12348 13277 12357 13311
rect 12357 13277 12391 13311
rect 12391 13277 12400 13311
rect 12348 13268 12400 13277
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 13636 13268 13688 13320
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 10784 13243 10836 13252
rect 10784 13209 10793 13243
rect 10793 13209 10827 13243
rect 10827 13209 10836 13243
rect 10784 13200 10836 13209
rect 12072 13200 12124 13252
rect 3516 13132 3568 13184
rect 7288 13132 7340 13184
rect 11520 13132 11572 13184
rect 12900 13175 12952 13184
rect 12900 13141 12909 13175
rect 12909 13141 12943 13175
rect 12943 13141 12952 13175
rect 12900 13132 12952 13141
rect 15384 13200 15436 13252
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 18880 13404 18932 13456
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 17868 13336 17920 13388
rect 19800 13472 19852 13524
rect 20352 13515 20404 13524
rect 20352 13481 20361 13515
rect 20361 13481 20395 13515
rect 20395 13481 20404 13515
rect 20352 13472 20404 13481
rect 25044 13472 25096 13524
rect 19432 13404 19484 13456
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 17960 13200 18012 13252
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 18788 13311 18840 13320
rect 18788 13277 18797 13311
rect 18797 13277 18831 13311
rect 18831 13277 18840 13311
rect 18788 13268 18840 13277
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 15200 13132 15252 13184
rect 17132 13132 17184 13184
rect 17592 13132 17644 13184
rect 18052 13132 18104 13184
rect 18604 13132 18656 13184
rect 19064 13268 19116 13320
rect 20168 13268 20220 13320
rect 20720 13336 20772 13388
rect 25780 13311 25832 13320
rect 25780 13277 25789 13311
rect 25789 13277 25823 13311
rect 25823 13277 25832 13311
rect 25780 13268 25832 13277
rect 21088 13243 21140 13252
rect 21088 13209 21097 13243
rect 21097 13209 21131 13243
rect 21131 13209 21140 13243
rect 21088 13200 21140 13209
rect 23112 13200 23164 13252
rect 22376 13132 22428 13184
rect 4761 13030 4813 13082
rect 4825 13030 4877 13082
rect 4889 13030 4941 13082
rect 4953 13030 5005 13082
rect 5017 13030 5069 13082
rect 11063 13030 11115 13082
rect 11127 13030 11179 13082
rect 11191 13030 11243 13082
rect 11255 13030 11307 13082
rect 11319 13030 11371 13082
rect 17365 13030 17417 13082
rect 17429 13030 17481 13082
rect 17493 13030 17545 13082
rect 17557 13030 17609 13082
rect 17621 13030 17673 13082
rect 23667 13030 23719 13082
rect 23731 13030 23783 13082
rect 23795 13030 23847 13082
rect 23859 13030 23911 13082
rect 23923 13030 23975 13082
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 4436 12928 4488 12980
rect 4804 12928 4856 12980
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 2228 12792 2280 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 4436 12792 4488 12844
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 6552 12724 6604 12776
rect 5264 12656 5316 12708
rect 6736 12656 6788 12708
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 8576 12792 8628 12844
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 8392 12656 8444 12708
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 12808 12928 12860 12980
rect 13084 12928 13136 12980
rect 14280 12928 14332 12980
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 17776 12928 17828 12980
rect 17960 12928 18012 12980
rect 18236 12928 18288 12980
rect 18604 12971 18656 12980
rect 18604 12937 18613 12971
rect 18613 12937 18647 12971
rect 18647 12937 18656 12971
rect 18604 12928 18656 12937
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 23112 12971 23164 12980
rect 23112 12937 23121 12971
rect 23121 12937 23155 12971
rect 23155 12937 23164 12971
rect 23112 12928 23164 12937
rect 9956 12860 10008 12912
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 10140 12835 10192 12844
rect 10140 12801 10149 12835
rect 10149 12801 10183 12835
rect 10183 12801 10192 12835
rect 10140 12792 10192 12801
rect 8944 12724 8996 12776
rect 10876 12903 10928 12912
rect 10876 12869 10885 12903
rect 10885 12869 10919 12903
rect 10919 12869 10928 12903
rect 10876 12860 10928 12869
rect 12900 12860 12952 12912
rect 11060 12835 11112 12844
rect 11060 12801 11069 12835
rect 11069 12801 11103 12835
rect 11103 12801 11112 12835
rect 11060 12792 11112 12801
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 11888 12792 11940 12844
rect 15568 12792 15620 12844
rect 16028 12792 16080 12844
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 18052 12860 18104 12912
rect 18880 12792 18932 12844
rect 20352 12792 20404 12844
rect 21180 12792 21232 12844
rect 24676 12792 24728 12844
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 5540 12588 5592 12640
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 7472 12588 7524 12640
rect 8300 12588 8352 12640
rect 9680 12656 9732 12708
rect 9772 12656 9824 12708
rect 11704 12724 11756 12776
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 16488 12724 16540 12776
rect 16396 12656 16448 12708
rect 17224 12724 17276 12776
rect 18236 12724 18288 12776
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 21548 12767 21600 12776
rect 21548 12733 21557 12767
rect 21557 12733 21591 12767
rect 21591 12733 21600 12767
rect 21548 12724 21600 12733
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 11612 12588 11664 12640
rect 11796 12588 11848 12640
rect 18144 12656 18196 12708
rect 17776 12631 17828 12640
rect 17776 12597 17785 12631
rect 17785 12597 17819 12631
rect 17819 12597 17828 12631
rect 17776 12588 17828 12597
rect 22284 12588 22336 12640
rect 4101 12486 4153 12538
rect 4165 12486 4217 12538
rect 4229 12486 4281 12538
rect 4293 12486 4345 12538
rect 4357 12486 4409 12538
rect 10403 12486 10455 12538
rect 10467 12486 10519 12538
rect 10531 12486 10583 12538
rect 10595 12486 10647 12538
rect 10659 12486 10711 12538
rect 16705 12486 16757 12538
rect 16769 12486 16821 12538
rect 16833 12486 16885 12538
rect 16897 12486 16949 12538
rect 16961 12486 17013 12538
rect 23007 12486 23059 12538
rect 23071 12486 23123 12538
rect 23135 12486 23187 12538
rect 23199 12486 23251 12538
rect 23263 12486 23315 12538
rect 3056 12384 3108 12436
rect 3424 12384 3476 12436
rect 6184 12384 6236 12436
rect 7288 12384 7340 12436
rect 12164 12384 12216 12436
rect 13544 12384 13596 12436
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 17040 12384 17092 12436
rect 4804 12359 4856 12368
rect 4804 12325 4813 12359
rect 4813 12325 4847 12359
rect 4847 12325 4856 12359
rect 4804 12316 4856 12325
rect 2136 12291 2188 12300
rect 2136 12257 2145 12291
rect 2145 12257 2179 12291
rect 2179 12257 2188 12291
rect 2136 12248 2188 12257
rect 3516 12248 3568 12300
rect 3884 12180 3936 12232
rect 5540 12248 5592 12300
rect 8484 12359 8536 12368
rect 8484 12325 8493 12359
rect 8493 12325 8527 12359
rect 8527 12325 8536 12359
rect 8484 12316 8536 12325
rect 16396 12316 16448 12368
rect 17316 12316 17368 12368
rect 6552 12248 6604 12300
rect 8208 12248 8260 12300
rect 5172 12180 5224 12232
rect 5448 12180 5500 12232
rect 6092 12223 6144 12232
rect 6092 12189 6099 12223
rect 6099 12189 6144 12223
rect 6092 12180 6144 12189
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 2504 12112 2556 12164
rect 2688 12112 2740 12164
rect 4344 12112 4396 12164
rect 5816 12112 5868 12164
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 3792 12044 3844 12096
rect 5356 12044 5408 12096
rect 6000 12044 6052 12096
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 8300 12180 8352 12232
rect 8576 12180 8628 12232
rect 11520 12248 11572 12300
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 11612 12180 11664 12232
rect 9220 12112 9272 12164
rect 11888 12180 11940 12232
rect 16028 12180 16080 12232
rect 21364 12248 21416 12300
rect 22468 12248 22520 12300
rect 13176 12112 13228 12164
rect 17776 12180 17828 12232
rect 20720 12223 20772 12232
rect 20720 12189 20729 12223
rect 20729 12189 20763 12223
rect 20763 12189 20772 12223
rect 20720 12180 20772 12189
rect 24676 12180 24728 12232
rect 18236 12112 18288 12164
rect 20904 12112 20956 12164
rect 22284 12112 22336 12164
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 7656 12044 7708 12096
rect 9588 12044 9640 12096
rect 14556 12044 14608 12096
rect 21180 12044 21232 12096
rect 21916 12044 21968 12096
rect 22008 12044 22060 12096
rect 24492 12087 24544 12096
rect 24492 12053 24501 12087
rect 24501 12053 24535 12087
rect 24535 12053 24544 12087
rect 24492 12044 24544 12053
rect 4761 11942 4813 11994
rect 4825 11942 4877 11994
rect 4889 11942 4941 11994
rect 4953 11942 5005 11994
rect 5017 11942 5069 11994
rect 11063 11942 11115 11994
rect 11127 11942 11179 11994
rect 11191 11942 11243 11994
rect 11255 11942 11307 11994
rect 11319 11942 11371 11994
rect 17365 11942 17417 11994
rect 17429 11942 17481 11994
rect 17493 11942 17545 11994
rect 17557 11942 17609 11994
rect 17621 11942 17673 11994
rect 23667 11942 23719 11994
rect 23731 11942 23783 11994
rect 23795 11942 23847 11994
rect 23859 11942 23911 11994
rect 23923 11942 23975 11994
rect 2412 11840 2464 11892
rect 2044 11772 2096 11824
rect 2596 11704 2648 11756
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3240 11747 3292 11756
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 4344 11883 4396 11892
rect 4344 11849 4353 11883
rect 4353 11849 4387 11883
rect 4387 11849 4396 11883
rect 4344 11840 4396 11849
rect 5816 11883 5868 11892
rect 5816 11849 5825 11883
rect 5825 11849 5859 11883
rect 5859 11849 5868 11883
rect 5816 11840 5868 11849
rect 6092 11840 6144 11892
rect 6644 11840 6696 11892
rect 8392 11840 8444 11892
rect 10140 11840 10192 11892
rect 10784 11840 10836 11892
rect 11520 11840 11572 11892
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 3976 11772 4028 11824
rect 5540 11815 5592 11824
rect 5540 11781 5549 11815
rect 5549 11781 5583 11815
rect 5583 11781 5592 11815
rect 5540 11772 5592 11781
rect 6276 11772 6328 11824
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 4896 11704 4948 11756
rect 2228 11568 2280 11620
rect 2504 11611 2556 11620
rect 2504 11577 2513 11611
rect 2513 11577 2547 11611
rect 2547 11577 2556 11611
rect 2504 11568 2556 11577
rect 3884 11611 3936 11620
rect 3884 11577 3893 11611
rect 3893 11577 3927 11611
rect 3927 11577 3936 11611
rect 3884 11568 3936 11577
rect 4436 11568 4488 11620
rect 5637 11747 5689 11756
rect 5637 11713 5646 11747
rect 5646 11713 5680 11747
rect 5680 11713 5689 11747
rect 5637 11704 5689 11713
rect 6092 11704 6144 11756
rect 7380 11772 7432 11824
rect 8116 11772 8168 11824
rect 6736 11704 6788 11756
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 9588 11747 9640 11756
rect 9588 11713 9597 11747
rect 9597 11713 9631 11747
rect 9631 11713 9640 11747
rect 9588 11704 9640 11713
rect 6000 11636 6052 11688
rect 7196 11636 7248 11688
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 9220 11679 9272 11688
rect 9220 11645 9229 11679
rect 9229 11645 9263 11679
rect 9263 11645 9272 11679
rect 9220 11636 9272 11645
rect 10048 11636 10100 11688
rect 6276 11568 6328 11620
rect 10968 11568 11020 11620
rect 11980 11704 12032 11756
rect 12072 11704 12124 11756
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 14096 11704 14148 11756
rect 14832 11840 14884 11892
rect 14556 11815 14608 11824
rect 14556 11781 14565 11815
rect 14565 11781 14599 11815
rect 14599 11781 14608 11815
rect 14556 11772 14608 11781
rect 18788 11883 18840 11892
rect 18788 11849 18813 11883
rect 18813 11849 18840 11883
rect 18788 11840 18840 11849
rect 20904 11883 20956 11892
rect 20904 11849 20913 11883
rect 20913 11849 20947 11883
rect 20947 11849 20956 11883
rect 20904 11840 20956 11849
rect 17132 11772 17184 11824
rect 17776 11772 17828 11824
rect 18420 11772 18472 11824
rect 21456 11840 21508 11892
rect 21548 11840 21600 11892
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 12992 11636 13044 11688
rect 15568 11636 15620 11688
rect 20812 11704 20864 11756
rect 12164 11568 12216 11620
rect 15660 11568 15712 11620
rect 18328 11636 18380 11688
rect 21180 11747 21232 11756
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 20996 11636 21048 11688
rect 21364 11747 21416 11756
rect 21364 11713 21399 11747
rect 21399 11713 21416 11747
rect 21364 11704 21416 11713
rect 21916 11772 21968 11824
rect 23480 11840 23532 11892
rect 21824 11704 21876 11756
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 22192 11772 22244 11824
rect 24492 11772 24544 11824
rect 22376 11704 22428 11756
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 22928 11704 22980 11756
rect 23112 11747 23164 11756
rect 23112 11713 23121 11747
rect 23121 11713 23155 11747
rect 23155 11713 23164 11747
rect 23112 11704 23164 11713
rect 24584 11704 24636 11756
rect 5908 11500 5960 11552
rect 6736 11500 6788 11552
rect 11520 11500 11572 11552
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 18236 11500 18288 11552
rect 24032 11636 24084 11688
rect 21640 11568 21692 11620
rect 19432 11500 19484 11552
rect 20904 11500 20956 11552
rect 21456 11500 21508 11552
rect 21824 11500 21876 11552
rect 22008 11500 22060 11552
rect 23940 11500 23992 11552
rect 24952 11568 25004 11620
rect 25688 11543 25740 11552
rect 25688 11509 25697 11543
rect 25697 11509 25731 11543
rect 25731 11509 25740 11543
rect 25688 11500 25740 11509
rect 4101 11398 4153 11450
rect 4165 11398 4217 11450
rect 4229 11398 4281 11450
rect 4293 11398 4345 11450
rect 4357 11398 4409 11450
rect 10403 11398 10455 11450
rect 10467 11398 10519 11450
rect 10531 11398 10583 11450
rect 10595 11398 10647 11450
rect 10659 11398 10711 11450
rect 16705 11398 16757 11450
rect 16769 11398 16821 11450
rect 16833 11398 16885 11450
rect 16897 11398 16949 11450
rect 16961 11398 17013 11450
rect 23007 11398 23059 11450
rect 23071 11398 23123 11450
rect 23135 11398 23187 11450
rect 23199 11398 23251 11450
rect 23263 11398 23315 11450
rect 3056 11296 3108 11348
rect 4620 11296 4672 11348
rect 4896 11339 4948 11348
rect 4896 11305 4905 11339
rect 4905 11305 4939 11339
rect 4939 11305 4948 11339
rect 4896 11296 4948 11305
rect 3332 11228 3384 11280
rect 5264 11271 5316 11280
rect 5264 11237 5273 11271
rect 5273 11237 5307 11271
rect 5307 11237 5316 11271
rect 5264 11228 5316 11237
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 6276 11296 6328 11348
rect 8576 11296 8628 11348
rect 8852 11296 8904 11348
rect 5540 11228 5592 11280
rect 5724 11228 5776 11280
rect 6368 11271 6420 11280
rect 6368 11237 6377 11271
rect 6377 11237 6411 11271
rect 6411 11237 6420 11271
rect 6368 11228 6420 11237
rect 5172 11160 5224 11212
rect 6276 11160 6328 11212
rect 3240 11092 3292 11144
rect 6184 11092 6236 11144
rect 7196 11160 7248 11212
rect 9772 11160 9824 11212
rect 6552 11092 6604 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 6460 11024 6512 11076
rect 8484 11024 8536 11076
rect 9956 11024 10008 11076
rect 11060 11296 11112 11348
rect 11612 11339 11664 11348
rect 11612 11305 11621 11339
rect 11621 11305 11655 11339
rect 11655 11305 11664 11339
rect 11612 11296 11664 11305
rect 11796 11296 11848 11348
rect 11980 11228 12032 11280
rect 11704 11160 11756 11212
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 15660 11339 15712 11348
rect 10968 11092 11020 11144
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12440 11092 12492 11144
rect 11704 11024 11756 11076
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 16580 11228 16632 11280
rect 17776 11296 17828 11348
rect 13820 11092 13872 11144
rect 17960 11160 18012 11212
rect 18052 11160 18104 11212
rect 18328 11203 18380 11212
rect 18328 11169 18337 11203
rect 18337 11169 18371 11203
rect 18371 11169 18380 11203
rect 18328 11160 18380 11169
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 15568 11092 15620 11144
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20812 11296 20864 11348
rect 22284 11296 22336 11348
rect 21180 11228 21232 11280
rect 22008 11160 22060 11212
rect 22192 11160 22244 11212
rect 24032 11339 24084 11348
rect 23572 11228 23624 11280
rect 15476 11067 15528 11076
rect 15476 11033 15485 11067
rect 15485 11033 15519 11067
rect 15519 11033 15528 11067
rect 15476 11024 15528 11033
rect 4436 10956 4488 11008
rect 5264 10956 5316 11008
rect 6092 10956 6144 11008
rect 13636 10956 13688 11008
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 16028 11024 16080 11076
rect 17040 11024 17092 11076
rect 18696 11024 18748 11076
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 21548 11092 21600 11101
rect 18420 10956 18472 11008
rect 18788 10956 18840 11008
rect 21272 11024 21324 11076
rect 21824 11135 21876 11144
rect 21824 11101 21833 11135
rect 21833 11101 21867 11135
rect 21867 11101 21876 11135
rect 21824 11092 21876 11101
rect 23480 11160 23532 11212
rect 24032 11305 24041 11339
rect 24041 11305 24075 11339
rect 24075 11305 24084 11339
rect 24032 11296 24084 11305
rect 22928 11092 22980 11144
rect 21364 10956 21416 11008
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24032 11092 24084 11101
rect 24216 11135 24268 11144
rect 24216 11101 24225 11135
rect 24225 11101 24259 11135
rect 24259 11101 24268 11135
rect 24216 11092 24268 11101
rect 25688 11160 25740 11212
rect 24124 11024 24176 11076
rect 24216 10956 24268 11008
rect 4761 10854 4813 10906
rect 4825 10854 4877 10906
rect 4889 10854 4941 10906
rect 4953 10854 5005 10906
rect 5017 10854 5069 10906
rect 11063 10854 11115 10906
rect 11127 10854 11179 10906
rect 11191 10854 11243 10906
rect 11255 10854 11307 10906
rect 11319 10854 11371 10906
rect 17365 10854 17417 10906
rect 17429 10854 17481 10906
rect 17493 10854 17545 10906
rect 17557 10854 17609 10906
rect 17621 10854 17673 10906
rect 23667 10854 23719 10906
rect 23731 10854 23783 10906
rect 23795 10854 23847 10906
rect 23859 10854 23911 10906
rect 23923 10854 23975 10906
rect 5448 10752 5500 10804
rect 9312 10752 9364 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 17960 10752 18012 10804
rect 18328 10752 18380 10804
rect 2412 10727 2464 10736
rect 2412 10693 2421 10727
rect 2421 10693 2455 10727
rect 2455 10693 2464 10727
rect 2412 10684 2464 10693
rect 2872 10684 2924 10736
rect 6276 10684 6328 10736
rect 22192 10795 22244 10804
rect 22192 10761 22201 10795
rect 22201 10761 22235 10795
rect 22235 10761 22244 10795
rect 22192 10752 22244 10761
rect 24124 10752 24176 10804
rect 4528 10616 4580 10668
rect 4620 10616 4672 10668
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 5172 10480 5224 10532
rect 8576 10548 8628 10600
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9496 10616 9548 10668
rect 10876 10616 10928 10668
rect 9680 10548 9732 10600
rect 13636 10616 13688 10668
rect 14372 10616 14424 10668
rect 14924 10616 14976 10668
rect 15568 10616 15620 10668
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 15292 10548 15344 10600
rect 16304 10548 16356 10600
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 18972 10616 19024 10668
rect 19064 10659 19116 10668
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 2780 10412 2832 10421
rect 5356 10412 5408 10464
rect 5632 10412 5684 10464
rect 12808 10480 12860 10532
rect 13084 10480 13136 10532
rect 18604 10480 18656 10532
rect 19432 10548 19484 10600
rect 20996 10616 21048 10668
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 22284 10659 22336 10668
rect 22284 10625 22293 10659
rect 22293 10625 22327 10659
rect 22327 10625 22336 10659
rect 22284 10616 22336 10625
rect 23664 10659 23716 10668
rect 23664 10625 23673 10659
rect 23673 10625 23707 10659
rect 23707 10625 23716 10659
rect 23664 10616 23716 10625
rect 23848 10659 23900 10668
rect 23848 10625 23857 10659
rect 23857 10625 23891 10659
rect 23891 10625 23900 10659
rect 23848 10616 23900 10625
rect 23480 10548 23532 10600
rect 24216 10616 24268 10668
rect 24492 10659 24544 10668
rect 24492 10625 24501 10659
rect 24501 10625 24535 10659
rect 24535 10625 24544 10659
rect 24492 10616 24544 10625
rect 24768 10659 24820 10668
rect 24768 10625 24777 10659
rect 24777 10625 24811 10659
rect 24811 10625 24820 10659
rect 24768 10616 24820 10625
rect 24952 10659 25004 10668
rect 24952 10625 24961 10659
rect 24961 10625 24995 10659
rect 24995 10625 25004 10659
rect 24952 10616 25004 10625
rect 24584 10548 24636 10600
rect 13176 10412 13228 10464
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 15752 10412 15804 10464
rect 19708 10412 19760 10464
rect 21088 10412 21140 10464
rect 24124 10412 24176 10464
rect 4101 10310 4153 10362
rect 4165 10310 4217 10362
rect 4229 10310 4281 10362
rect 4293 10310 4345 10362
rect 4357 10310 4409 10362
rect 10403 10310 10455 10362
rect 10467 10310 10519 10362
rect 10531 10310 10583 10362
rect 10595 10310 10647 10362
rect 10659 10310 10711 10362
rect 16705 10310 16757 10362
rect 16769 10310 16821 10362
rect 16833 10310 16885 10362
rect 16897 10310 16949 10362
rect 16961 10310 17013 10362
rect 23007 10310 23059 10362
rect 23071 10310 23123 10362
rect 23135 10310 23187 10362
rect 23199 10310 23251 10362
rect 23263 10310 23315 10362
rect 6736 10208 6788 10260
rect 6920 10208 6972 10260
rect 8944 10208 8996 10260
rect 11980 10251 12032 10260
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 13544 10208 13596 10260
rect 14740 10208 14792 10260
rect 16948 10208 17000 10260
rect 18328 10208 18380 10260
rect 18604 10208 18656 10260
rect 2136 10140 2188 10192
rect 13728 10140 13780 10192
rect 15660 10140 15712 10192
rect 17040 10140 17092 10192
rect 12808 10072 12860 10124
rect 2780 10004 2832 10056
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 5908 10004 5960 10056
rect 6000 9936 6052 9988
rect 6828 9936 6880 9988
rect 3792 9868 3844 9920
rect 6368 9868 6420 9920
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 9128 10004 9180 10056
rect 9680 10004 9732 10056
rect 10968 10004 11020 10056
rect 11520 10004 11572 10056
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 13360 10072 13412 10124
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 13912 10072 13964 10124
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13636 10004 13688 10056
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 14464 10004 14516 10056
rect 14924 10004 14976 10056
rect 12808 9936 12860 9988
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 7564 9868 7616 9877
rect 13176 9868 13228 9920
rect 13360 9979 13412 9988
rect 13360 9945 13369 9979
rect 13369 9945 13403 9979
rect 13403 9945 13412 9979
rect 13360 9936 13412 9945
rect 13820 9936 13872 9988
rect 16396 10004 16448 10056
rect 16672 10047 16724 10056
rect 16672 10013 16681 10047
rect 16681 10013 16715 10047
rect 16715 10013 16724 10047
rect 16672 10004 16724 10013
rect 16304 9979 16356 9988
rect 16304 9945 16313 9979
rect 16313 9945 16347 9979
rect 16347 9945 16356 9979
rect 16304 9936 16356 9945
rect 18512 10140 18564 10192
rect 18144 9936 18196 9988
rect 19064 10004 19116 10056
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 17132 9868 17184 9920
rect 18052 9868 18104 9920
rect 19708 10004 19760 10056
rect 20904 10208 20956 10260
rect 21824 10208 21876 10260
rect 20720 10140 20772 10192
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 21088 10115 21140 10124
rect 21088 10081 21097 10115
rect 21097 10081 21131 10115
rect 21131 10081 21140 10115
rect 21088 10072 21140 10081
rect 22928 10208 22980 10260
rect 24492 10208 24544 10260
rect 24768 10208 24820 10260
rect 23848 10140 23900 10192
rect 20628 10004 20680 10056
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 23388 10047 23440 10056
rect 23388 10013 23397 10047
rect 23397 10013 23431 10047
rect 23431 10013 23440 10047
rect 23388 10004 23440 10013
rect 24492 10115 24544 10124
rect 24492 10081 24501 10115
rect 24501 10081 24535 10115
rect 24535 10081 24544 10115
rect 24492 10072 24544 10081
rect 24676 10072 24728 10124
rect 24860 10004 24912 10056
rect 25136 10004 25188 10056
rect 20996 9936 21048 9988
rect 22376 9936 22428 9988
rect 21364 9868 21416 9920
rect 22560 9911 22612 9920
rect 22560 9877 22569 9911
rect 22569 9877 22603 9911
rect 22603 9877 22612 9911
rect 23664 9936 23716 9988
rect 24492 9936 24544 9988
rect 22560 9868 22612 9877
rect 23296 9868 23348 9920
rect 25412 9911 25464 9920
rect 25412 9877 25421 9911
rect 25421 9877 25455 9911
rect 25455 9877 25464 9911
rect 25412 9868 25464 9877
rect 4761 9766 4813 9818
rect 4825 9766 4877 9818
rect 4889 9766 4941 9818
rect 4953 9766 5005 9818
rect 5017 9766 5069 9818
rect 11063 9766 11115 9818
rect 11127 9766 11179 9818
rect 11191 9766 11243 9818
rect 11255 9766 11307 9818
rect 11319 9766 11371 9818
rect 17365 9766 17417 9818
rect 17429 9766 17481 9818
rect 17493 9766 17545 9818
rect 17557 9766 17609 9818
rect 17621 9766 17673 9818
rect 23667 9766 23719 9818
rect 23731 9766 23783 9818
rect 23795 9766 23847 9818
rect 23859 9766 23911 9818
rect 23923 9766 23975 9818
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 2136 9528 2188 9580
rect 2320 9528 2372 9580
rect 3792 9528 3844 9580
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 5632 9596 5684 9648
rect 6000 9639 6052 9648
rect 6000 9605 6009 9639
rect 6009 9605 6043 9639
rect 6043 9605 6052 9639
rect 6000 9596 6052 9605
rect 6552 9664 6604 9716
rect 13360 9664 13412 9716
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 3516 9460 3568 9512
rect 6092 9528 6144 9580
rect 7564 9528 7616 9580
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 8024 9528 8076 9537
rect 2504 9324 2556 9376
rect 3424 9324 3476 9376
rect 4436 9324 4488 9376
rect 5080 9324 5132 9376
rect 5448 9460 5500 9512
rect 9496 9528 9548 9580
rect 10876 9528 10928 9580
rect 11704 9596 11756 9648
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 13176 9596 13228 9648
rect 12164 9528 12216 9580
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 15384 9596 15436 9648
rect 16120 9596 16172 9648
rect 10968 9460 11020 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 12900 9392 12952 9444
rect 5816 9324 5868 9376
rect 6276 9324 6328 9376
rect 10324 9324 10376 9376
rect 12348 9324 12400 9376
rect 13176 9367 13228 9376
rect 13176 9333 13185 9367
rect 13185 9333 13219 9367
rect 13219 9333 13228 9367
rect 13176 9324 13228 9333
rect 13820 9392 13872 9444
rect 14096 9528 14148 9580
rect 14372 9528 14424 9580
rect 14924 9571 14976 9580
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 16212 9528 16264 9580
rect 16672 9596 16724 9648
rect 16304 9460 16356 9512
rect 14188 9392 14240 9444
rect 16396 9392 16448 9444
rect 17224 9596 17276 9648
rect 18236 9664 18288 9716
rect 18604 9596 18656 9648
rect 18696 9639 18748 9648
rect 18696 9605 18705 9639
rect 18705 9605 18739 9639
rect 18739 9605 18748 9639
rect 18696 9596 18748 9605
rect 18144 9528 18196 9580
rect 18880 9571 18932 9580
rect 18880 9537 18889 9571
rect 18889 9537 18923 9571
rect 18923 9537 18932 9571
rect 18880 9528 18932 9537
rect 20628 9596 20680 9648
rect 20720 9639 20772 9648
rect 20720 9605 20729 9639
rect 20729 9605 20763 9639
rect 20763 9605 20772 9639
rect 22100 9664 22152 9716
rect 23388 9664 23440 9716
rect 20720 9596 20772 9605
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 19340 9571 19392 9580
rect 19340 9537 19349 9571
rect 19349 9537 19383 9571
rect 19383 9537 19392 9571
rect 19340 9528 19392 9537
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 16948 9392 17000 9444
rect 15292 9367 15344 9376
rect 15292 9333 15301 9367
rect 15301 9333 15335 9367
rect 15335 9333 15344 9367
rect 15292 9324 15344 9333
rect 17868 9392 17920 9444
rect 18696 9392 18748 9444
rect 20720 9392 20772 9444
rect 21364 9571 21416 9580
rect 21364 9537 21373 9571
rect 21373 9537 21407 9571
rect 21407 9537 21416 9571
rect 21364 9528 21416 9537
rect 21548 9571 21600 9580
rect 21548 9537 21557 9571
rect 21557 9537 21591 9571
rect 21591 9537 21600 9571
rect 21548 9528 21600 9537
rect 21824 9528 21876 9580
rect 22100 9571 22152 9580
rect 22100 9537 22109 9571
rect 22109 9537 22143 9571
rect 22143 9537 22152 9571
rect 22100 9528 22152 9537
rect 24124 9596 24176 9648
rect 25412 9596 25464 9648
rect 22560 9528 22612 9580
rect 21456 9503 21508 9512
rect 21456 9469 21465 9503
rect 21465 9469 21499 9503
rect 21499 9469 21508 9503
rect 21456 9460 21508 9469
rect 23388 9460 23440 9512
rect 24860 9460 24912 9512
rect 22468 9392 22520 9444
rect 23296 9392 23348 9444
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 17684 9324 17736 9376
rect 18328 9324 18380 9376
rect 18420 9367 18472 9376
rect 18420 9333 18429 9367
rect 18429 9333 18463 9367
rect 18463 9333 18472 9367
rect 18420 9324 18472 9333
rect 18880 9324 18932 9376
rect 19616 9324 19668 9376
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 21548 9324 21600 9376
rect 22284 9324 22336 9376
rect 23480 9324 23532 9376
rect 25136 9324 25188 9376
rect 4101 9222 4153 9274
rect 4165 9222 4217 9274
rect 4229 9222 4281 9274
rect 4293 9222 4345 9274
rect 4357 9222 4409 9274
rect 10403 9222 10455 9274
rect 10467 9222 10519 9274
rect 10531 9222 10583 9274
rect 10595 9222 10647 9274
rect 10659 9222 10711 9274
rect 16705 9222 16757 9274
rect 16769 9222 16821 9274
rect 16833 9222 16885 9274
rect 16897 9222 16949 9274
rect 16961 9222 17013 9274
rect 23007 9222 23059 9274
rect 23071 9222 23123 9274
rect 23135 9222 23187 9274
rect 23199 9222 23251 9274
rect 23263 9222 23315 9274
rect 2320 9120 2372 9172
rect 2596 9120 2648 9172
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3516 9163 3568 9172
rect 1768 9052 1820 9104
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 4620 9120 4672 9172
rect 4160 9095 4212 9104
rect 4160 9061 4169 9095
rect 4169 9061 4203 9095
rect 4203 9061 4212 9095
rect 4160 9052 4212 9061
rect 4436 9052 4488 9104
rect 4804 9095 4856 9104
rect 4804 9061 4813 9095
rect 4813 9061 4847 9095
rect 4847 9061 4856 9095
rect 4804 9052 4856 9061
rect 1860 8984 1912 9036
rect 2688 8984 2740 9036
rect 2320 8891 2372 8900
rect 2320 8857 2329 8891
rect 2329 8857 2363 8891
rect 2363 8857 2372 8891
rect 2320 8848 2372 8857
rect 2504 8891 2556 8900
rect 2504 8857 2529 8891
rect 2529 8857 2556 8891
rect 2504 8848 2556 8857
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 4620 8916 4672 8968
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 8024 9120 8076 9172
rect 11520 9120 11572 9172
rect 11888 9120 11940 9172
rect 12808 9120 12860 9172
rect 12992 9120 13044 9172
rect 13176 9120 13228 9172
rect 13268 9120 13320 9172
rect 14004 9120 14056 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 5632 9052 5684 9104
rect 5908 8984 5960 9036
rect 6000 9027 6052 9036
rect 6000 8993 6009 9027
rect 6009 8993 6043 9027
rect 6043 8993 6052 9027
rect 6000 8984 6052 8993
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 5724 8959 5776 8964
rect 3792 8891 3844 8900
rect 3792 8857 3801 8891
rect 3801 8857 3835 8891
rect 3835 8857 3844 8891
rect 3792 8848 3844 8857
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 5724 8925 5750 8959
rect 5750 8925 5776 8959
rect 5724 8912 5776 8925
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6460 8984 6512 9036
rect 8116 8984 8168 9036
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 6000 8848 6052 8900
rect 6552 8848 6604 8900
rect 9128 8916 9180 8968
rect 12440 8984 12492 9036
rect 11704 8916 11756 8968
rect 12256 8959 12308 8968
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 13452 9052 13504 9104
rect 13636 9052 13688 9104
rect 14188 9052 14240 9104
rect 12808 8984 12860 9036
rect 6736 8848 6788 8900
rect 10140 8891 10192 8900
rect 10140 8857 10174 8891
rect 10174 8857 10192 8891
rect 10140 8848 10192 8857
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 13084 8984 13136 9036
rect 13268 8984 13320 9036
rect 16396 9120 16448 9172
rect 17132 9120 17184 9172
rect 17500 9120 17552 9172
rect 18420 9120 18472 9172
rect 19340 9120 19392 9172
rect 20996 9120 21048 9172
rect 22100 9120 22152 9172
rect 19708 9052 19760 9104
rect 22376 9120 22428 9172
rect 22468 9052 22520 9104
rect 14832 9027 14884 9036
rect 14832 8993 14841 9027
rect 14841 8993 14875 9027
rect 14875 8993 14884 9027
rect 14832 8984 14884 8993
rect 16580 8984 16632 9036
rect 20812 8984 20864 9036
rect 6276 8780 6328 8832
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 14004 8916 14056 8968
rect 13084 8848 13136 8900
rect 13452 8848 13504 8900
rect 15200 8959 15252 8968
rect 15200 8925 15209 8959
rect 15209 8925 15243 8959
rect 15243 8925 15252 8959
rect 15200 8916 15252 8925
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 18696 8916 18748 8968
rect 19064 8916 19116 8968
rect 15752 8848 15804 8900
rect 13360 8780 13412 8832
rect 19156 8848 19208 8900
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 22560 8916 22612 8968
rect 24676 8916 24728 8968
rect 22652 8848 22704 8900
rect 16488 8780 16540 8832
rect 17868 8780 17920 8832
rect 18144 8780 18196 8832
rect 19340 8823 19392 8832
rect 19340 8789 19349 8823
rect 19349 8789 19383 8823
rect 19383 8789 19392 8823
rect 19340 8780 19392 8789
rect 24400 8780 24452 8832
rect 4761 8678 4813 8730
rect 4825 8678 4877 8730
rect 4889 8678 4941 8730
rect 4953 8678 5005 8730
rect 5017 8678 5069 8730
rect 11063 8678 11115 8730
rect 11127 8678 11179 8730
rect 11191 8678 11243 8730
rect 11255 8678 11307 8730
rect 11319 8678 11371 8730
rect 17365 8678 17417 8730
rect 17429 8678 17481 8730
rect 17493 8678 17545 8730
rect 17557 8678 17609 8730
rect 17621 8678 17673 8730
rect 23667 8678 23719 8730
rect 23731 8678 23783 8730
rect 23795 8678 23847 8730
rect 23859 8678 23911 8730
rect 23923 8678 23975 8730
rect 1952 8576 2004 8628
rect 4160 8576 4212 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 3240 8440 3292 8492
rect 4528 8508 4580 8560
rect 4620 8508 4672 8560
rect 4988 8576 5040 8628
rect 5448 8576 5500 8628
rect 5724 8576 5776 8628
rect 6920 8576 6972 8628
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 13452 8576 13504 8628
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 16396 8576 16448 8628
rect 20260 8576 20312 8628
rect 22652 8619 22704 8628
rect 22652 8585 22661 8619
rect 22661 8585 22695 8619
rect 22695 8585 22704 8619
rect 22652 8576 22704 8585
rect 25136 8619 25188 8628
rect 25136 8585 25145 8619
rect 25145 8585 25179 8619
rect 25179 8585 25188 8619
rect 25136 8576 25188 8585
rect 6276 8508 6328 8560
rect 11980 8508 12032 8560
rect 2320 8372 2372 8424
rect 2688 8304 2740 8356
rect 4712 8304 4764 8356
rect 2596 8236 2648 8288
rect 4620 8236 4672 8288
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 8392 8483 8444 8492
rect 8392 8449 8426 8483
rect 8426 8449 8444 8483
rect 8392 8440 8444 8449
rect 10876 8440 10928 8492
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12440 8508 12492 8560
rect 12808 8508 12860 8560
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13360 8440 13412 8492
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 14372 8508 14424 8560
rect 16488 8508 16540 8560
rect 16672 8551 16724 8560
rect 16672 8517 16681 8551
rect 16681 8517 16715 8551
rect 16715 8517 16724 8551
rect 16672 8508 16724 8517
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 15292 8440 15344 8492
rect 16212 8440 16264 8492
rect 18512 8508 18564 8560
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18328 8440 18380 8492
rect 20812 8508 20864 8560
rect 23572 8508 23624 8560
rect 24400 8508 24452 8560
rect 18788 8440 18840 8492
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 23388 8483 23440 8492
rect 23388 8449 23397 8483
rect 23397 8449 23431 8483
rect 23431 8449 23440 8483
rect 23388 8440 23440 8449
rect 5816 8304 5868 8356
rect 6828 8304 6880 8356
rect 12440 8304 12492 8356
rect 11888 8236 11940 8288
rect 12256 8236 12308 8288
rect 18052 8304 18104 8356
rect 19156 8304 19208 8356
rect 22468 8304 22520 8356
rect 25872 8347 25924 8356
rect 25872 8313 25881 8347
rect 25881 8313 25915 8347
rect 25915 8313 25924 8347
rect 25872 8304 25924 8313
rect 13268 8236 13320 8288
rect 14556 8236 14608 8288
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 16212 8236 16264 8288
rect 17132 8279 17184 8288
rect 17132 8245 17141 8279
rect 17141 8245 17175 8279
rect 17175 8245 17184 8279
rect 17132 8236 17184 8245
rect 18328 8279 18380 8288
rect 18328 8245 18337 8279
rect 18337 8245 18371 8279
rect 18371 8245 18380 8279
rect 18328 8236 18380 8245
rect 4101 8134 4153 8186
rect 4165 8134 4217 8186
rect 4229 8134 4281 8186
rect 4293 8134 4345 8186
rect 4357 8134 4409 8186
rect 10403 8134 10455 8186
rect 10467 8134 10519 8186
rect 10531 8134 10583 8186
rect 10595 8134 10647 8186
rect 10659 8134 10711 8186
rect 16705 8134 16757 8186
rect 16769 8134 16821 8186
rect 16833 8134 16885 8186
rect 16897 8134 16949 8186
rect 16961 8134 17013 8186
rect 23007 8134 23059 8186
rect 23071 8134 23123 8186
rect 23135 8134 23187 8186
rect 23199 8134 23251 8186
rect 23263 8134 23315 8186
rect 2596 8032 2648 8084
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 4712 8007 4764 8016
rect 4712 7973 4721 8007
rect 4721 7973 4755 8007
rect 4755 7973 4764 8007
rect 4712 7964 4764 7973
rect 3240 7803 3292 7812
rect 3240 7769 3249 7803
rect 3249 7769 3283 7803
rect 3283 7769 3292 7803
rect 3240 7760 3292 7769
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4252 7871 4304 7880
rect 4252 7837 4261 7871
rect 4261 7837 4295 7871
rect 4295 7837 4304 7871
rect 4252 7828 4304 7837
rect 4436 7760 4488 7812
rect 5172 7828 5224 7880
rect 5632 8007 5684 8016
rect 5632 7973 5641 8007
rect 5641 7973 5675 8007
rect 5675 7973 5684 8007
rect 6276 8075 6328 8084
rect 6276 8041 6285 8075
rect 6285 8041 6319 8075
rect 6319 8041 6328 8075
rect 6276 8032 6328 8041
rect 8392 8032 8444 8084
rect 10140 8032 10192 8084
rect 12900 8032 12952 8084
rect 5632 7964 5684 7973
rect 6368 7964 6420 8016
rect 5908 7896 5960 7948
rect 7656 7828 7708 7880
rect 9220 7828 9272 7880
rect 10232 7964 10284 8016
rect 10140 7896 10192 7948
rect 13912 8075 13964 8084
rect 13912 8041 13921 8075
rect 13921 8041 13955 8075
rect 13955 8041 13964 8075
rect 13912 8032 13964 8041
rect 15476 8032 15528 8084
rect 16212 8032 16264 8084
rect 16580 8032 16632 8084
rect 16488 7964 16540 8016
rect 18052 8075 18104 8084
rect 18052 8041 18061 8075
rect 18061 8041 18095 8075
rect 18095 8041 18104 8075
rect 18052 8032 18104 8041
rect 18420 8032 18472 8084
rect 19708 8075 19760 8084
rect 19708 8041 19717 8075
rect 19717 8041 19751 8075
rect 19751 8041 19760 8075
rect 19708 8032 19760 8041
rect 18144 7964 18196 8016
rect 18236 7964 18288 8016
rect 19524 8007 19576 8016
rect 19524 7973 19533 8007
rect 19533 7973 19567 8007
rect 19567 7973 19576 8007
rect 19524 7964 19576 7973
rect 12440 7828 12492 7880
rect 19340 7896 19392 7948
rect 5080 7760 5132 7812
rect 10048 7760 10100 7812
rect 3608 7735 3660 7744
rect 3608 7701 3617 7735
rect 3617 7701 3651 7735
rect 3651 7701 3660 7735
rect 3608 7692 3660 7701
rect 9864 7735 9916 7744
rect 9864 7701 9873 7735
rect 9873 7701 9907 7735
rect 9907 7701 9916 7735
rect 11796 7760 11848 7812
rect 9864 7692 9916 7701
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 17132 7828 17184 7880
rect 15660 7803 15712 7812
rect 15660 7769 15669 7803
rect 15669 7769 15703 7803
rect 15703 7769 15712 7803
rect 15660 7760 15712 7769
rect 17868 7828 17920 7880
rect 22652 7871 22704 7880
rect 22652 7837 22661 7871
rect 22661 7837 22695 7871
rect 22695 7837 22704 7871
rect 22652 7828 22704 7837
rect 15476 7692 15528 7744
rect 15568 7692 15620 7744
rect 17684 7760 17736 7812
rect 18420 7760 18472 7812
rect 18972 7760 19024 7812
rect 17868 7735 17920 7744
rect 17868 7701 17877 7735
rect 17877 7701 17911 7735
rect 17911 7701 17920 7735
rect 17868 7692 17920 7701
rect 17960 7692 18012 7744
rect 21456 7692 21508 7744
rect 4761 7590 4813 7642
rect 4825 7590 4877 7642
rect 4889 7590 4941 7642
rect 4953 7590 5005 7642
rect 5017 7590 5069 7642
rect 11063 7590 11115 7642
rect 11127 7590 11179 7642
rect 11191 7590 11243 7642
rect 11255 7590 11307 7642
rect 11319 7590 11371 7642
rect 17365 7590 17417 7642
rect 17429 7590 17481 7642
rect 17493 7590 17545 7642
rect 17557 7590 17609 7642
rect 17621 7590 17673 7642
rect 23667 7590 23719 7642
rect 23731 7590 23783 7642
rect 23795 7590 23847 7642
rect 23859 7590 23911 7642
rect 23923 7590 23975 7642
rect 4436 7488 4488 7540
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 10232 7488 10284 7540
rect 11796 7488 11848 7540
rect 18328 7488 18380 7540
rect 19156 7531 19208 7540
rect 19156 7497 19165 7531
rect 19165 7497 19199 7531
rect 19199 7497 19208 7531
rect 19156 7488 19208 7497
rect 10140 7420 10192 7472
rect 3608 7352 3660 7404
rect 4160 7352 4212 7404
rect 4620 7352 4672 7404
rect 8116 7352 8168 7404
rect 8944 7352 8996 7404
rect 12256 7420 12308 7472
rect 15292 7420 15344 7472
rect 16304 7420 16356 7472
rect 18420 7463 18472 7472
rect 18420 7429 18429 7463
rect 18429 7429 18463 7463
rect 18463 7429 18472 7463
rect 18420 7420 18472 7429
rect 18512 7420 18564 7472
rect 19800 7420 19852 7472
rect 22652 7488 22704 7540
rect 4344 7327 4396 7336
rect 4344 7293 4353 7327
rect 4353 7293 4387 7327
rect 4387 7293 4396 7327
rect 4344 7284 4396 7293
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 12440 7352 12492 7404
rect 12716 7352 12768 7404
rect 17868 7352 17920 7404
rect 22560 7420 22612 7472
rect 24032 7463 24084 7472
rect 24032 7429 24041 7463
rect 24041 7429 24075 7463
rect 24075 7429 24084 7463
rect 24032 7420 24084 7429
rect 24676 7420 24728 7472
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 21916 7352 21968 7404
rect 24308 7352 24360 7404
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 19340 7284 19392 7336
rect 19524 7284 19576 7336
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 20812 7327 20864 7336
rect 20812 7293 20821 7327
rect 20821 7293 20855 7327
rect 20855 7293 20864 7327
rect 20812 7284 20864 7293
rect 4528 7216 4580 7268
rect 9772 7216 9824 7268
rect 3792 7148 3844 7200
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 7472 7148 7524 7200
rect 9220 7148 9272 7200
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 19064 7259 19116 7268
rect 19064 7225 19073 7259
rect 19073 7225 19107 7259
rect 19107 7225 19116 7259
rect 19064 7216 19116 7225
rect 11152 7148 11204 7200
rect 11520 7148 11572 7200
rect 16120 7148 16172 7200
rect 17960 7148 18012 7200
rect 18236 7148 18288 7200
rect 18512 7148 18564 7200
rect 21272 7148 21324 7200
rect 4101 7046 4153 7098
rect 4165 7046 4217 7098
rect 4229 7046 4281 7098
rect 4293 7046 4345 7098
rect 4357 7046 4409 7098
rect 10403 7046 10455 7098
rect 10467 7046 10519 7098
rect 10531 7046 10583 7098
rect 10595 7046 10647 7098
rect 10659 7046 10711 7098
rect 16705 7046 16757 7098
rect 16769 7046 16821 7098
rect 16833 7046 16885 7098
rect 16897 7046 16949 7098
rect 16961 7046 17013 7098
rect 23007 7046 23059 7098
rect 23071 7046 23123 7098
rect 23135 7046 23187 7098
rect 23199 7046 23251 7098
rect 23263 7046 23315 7098
rect 5172 6987 5224 6996
rect 5172 6953 5181 6987
rect 5181 6953 5215 6987
rect 5215 6953 5224 6987
rect 5172 6944 5224 6953
rect 5448 6944 5500 6996
rect 6368 6944 6420 6996
rect 7380 6944 7432 6996
rect 7472 6987 7524 6996
rect 7472 6953 7481 6987
rect 7481 6953 7515 6987
rect 7515 6953 7524 6987
rect 7472 6944 7524 6953
rect 7656 6987 7708 6996
rect 7656 6953 7665 6987
rect 7665 6953 7699 6987
rect 7699 6953 7708 6987
rect 7656 6944 7708 6953
rect 9772 6944 9824 6996
rect 10968 6944 11020 6996
rect 7012 6808 7064 6860
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 10324 6808 10376 6860
rect 12256 6944 12308 6996
rect 15108 6944 15160 6996
rect 15384 6944 15436 6996
rect 15844 6944 15896 6996
rect 16212 6944 16264 6996
rect 16120 6876 16172 6928
rect 18420 6944 18472 6996
rect 19248 6944 19300 6996
rect 20536 6944 20588 6996
rect 20812 6944 20864 6996
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 5540 6740 5592 6792
rect 4712 6672 4764 6724
rect 7104 6740 7156 6792
rect 12900 6808 12952 6860
rect 17776 6808 17828 6860
rect 21916 6808 21968 6860
rect 22560 6808 22612 6860
rect 7196 6672 7248 6724
rect 9312 6672 9364 6724
rect 10968 6715 11020 6724
rect 10968 6681 10977 6715
rect 10977 6681 11011 6715
rect 11011 6681 11020 6715
rect 10968 6672 11020 6681
rect 12164 6672 12216 6724
rect 12716 6740 12768 6792
rect 12900 6672 12952 6724
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 15292 6740 15344 6792
rect 15752 6740 15804 6792
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 15568 6672 15620 6724
rect 16488 6672 16540 6724
rect 6552 6604 6604 6656
rect 6920 6604 6972 6656
rect 7840 6604 7892 6656
rect 9404 6604 9456 6656
rect 9680 6604 9732 6656
rect 11888 6604 11940 6656
rect 11980 6604 12032 6656
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 13268 6604 13320 6656
rect 15016 6604 15068 6656
rect 15476 6604 15528 6656
rect 18144 6740 18196 6792
rect 17868 6672 17920 6724
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 19708 6783 19760 6792
rect 19708 6749 19717 6783
rect 19717 6749 19751 6783
rect 19751 6749 19760 6783
rect 19708 6740 19760 6749
rect 21180 6740 21232 6792
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 19248 6604 19300 6656
rect 19800 6604 19852 6656
rect 23572 6604 23624 6656
rect 24124 6647 24176 6656
rect 24124 6613 24133 6647
rect 24133 6613 24167 6647
rect 24167 6613 24176 6647
rect 24124 6604 24176 6613
rect 4761 6502 4813 6554
rect 4825 6502 4877 6554
rect 4889 6502 4941 6554
rect 4953 6502 5005 6554
rect 5017 6502 5069 6554
rect 11063 6502 11115 6554
rect 11127 6502 11179 6554
rect 11191 6502 11243 6554
rect 11255 6502 11307 6554
rect 11319 6502 11371 6554
rect 17365 6502 17417 6554
rect 17429 6502 17481 6554
rect 17493 6502 17545 6554
rect 17557 6502 17609 6554
rect 17621 6502 17673 6554
rect 23667 6502 23719 6554
rect 23731 6502 23783 6554
rect 23795 6502 23847 6554
rect 23859 6502 23911 6554
rect 23923 6502 23975 6554
rect 5540 6400 5592 6452
rect 6644 6400 6696 6452
rect 6828 6400 6880 6452
rect 7656 6332 7708 6384
rect 5724 6307 5776 6316
rect 5724 6273 5731 6307
rect 5731 6273 5776 6307
rect 5724 6264 5776 6273
rect 6092 6264 6144 6316
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6828 6264 6880 6316
rect 5356 6171 5408 6180
rect 5356 6137 5365 6171
rect 5365 6137 5399 6171
rect 5399 6137 5408 6171
rect 5356 6128 5408 6137
rect 5632 6128 5684 6180
rect 6184 6171 6236 6180
rect 6184 6137 6193 6171
rect 6193 6137 6227 6171
rect 6227 6137 6236 6171
rect 6184 6128 6236 6137
rect 7288 6196 7340 6248
rect 8944 6443 8996 6452
rect 8944 6409 8953 6443
rect 8953 6409 8987 6443
rect 8987 6409 8996 6443
rect 8944 6400 8996 6409
rect 9220 6400 9272 6452
rect 9312 6400 9364 6452
rect 9864 6400 9916 6452
rect 10140 6400 10192 6452
rect 10232 6400 10284 6452
rect 11980 6400 12032 6452
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 15936 6400 15988 6452
rect 8300 6264 8352 6316
rect 9312 6264 9364 6316
rect 9404 6264 9456 6316
rect 7380 6171 7432 6180
rect 7380 6137 7389 6171
rect 7389 6137 7423 6171
rect 7423 6137 7432 6171
rect 7380 6128 7432 6137
rect 7564 6060 7616 6112
rect 8576 6128 8628 6180
rect 9680 6128 9732 6180
rect 8760 6060 8812 6112
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 10232 6264 10284 6316
rect 12256 6375 12308 6384
rect 12256 6341 12265 6375
rect 12265 6341 12299 6375
rect 12299 6341 12308 6375
rect 12256 6332 12308 6341
rect 12716 6375 12768 6384
rect 12716 6341 12725 6375
rect 12725 6341 12759 6375
rect 12759 6341 12768 6375
rect 12716 6332 12768 6341
rect 14188 6332 14240 6384
rect 14740 6332 14792 6384
rect 16120 6400 16172 6452
rect 17868 6400 17920 6452
rect 19340 6400 19392 6452
rect 19524 6400 19576 6452
rect 19708 6400 19760 6452
rect 10968 6264 11020 6316
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 15016 6264 15068 6316
rect 10324 6196 10376 6248
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 11060 6196 11112 6248
rect 11612 6196 11664 6248
rect 10048 6128 10100 6180
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 15936 6264 15988 6316
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 16304 6307 16356 6316
rect 16304 6273 16314 6307
rect 16314 6273 16348 6307
rect 16348 6273 16356 6307
rect 16304 6264 16356 6273
rect 16948 6264 17000 6316
rect 17224 6264 17276 6316
rect 18144 6264 18196 6316
rect 19248 6307 19300 6316
rect 19248 6273 19257 6307
rect 19257 6273 19291 6307
rect 19291 6273 19300 6307
rect 19248 6264 19300 6273
rect 19984 6332 20036 6384
rect 19524 6307 19576 6316
rect 19524 6273 19533 6307
rect 19533 6273 19567 6307
rect 19567 6273 19576 6307
rect 19524 6264 19576 6273
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 15292 6239 15344 6248
rect 15292 6205 15301 6239
rect 15301 6205 15335 6239
rect 15335 6205 15344 6239
rect 15292 6196 15344 6205
rect 15844 6196 15896 6248
rect 17040 6239 17092 6248
rect 17040 6205 17049 6239
rect 17049 6205 17083 6239
rect 17083 6205 17092 6239
rect 17040 6196 17092 6205
rect 19064 6196 19116 6248
rect 11336 6060 11388 6112
rect 14372 6060 14424 6112
rect 15108 6060 15160 6112
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 15936 6060 15988 6112
rect 17960 6128 18012 6180
rect 19340 6171 19392 6180
rect 19340 6137 19349 6171
rect 19349 6137 19383 6171
rect 19383 6137 19392 6171
rect 19340 6128 19392 6137
rect 20168 6307 20220 6316
rect 20168 6273 20177 6307
rect 20177 6273 20211 6307
rect 20211 6273 20220 6307
rect 20168 6264 20220 6273
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 20352 6196 20404 6248
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 20628 6196 20680 6248
rect 21272 6307 21324 6316
rect 21272 6273 21281 6307
rect 21281 6273 21315 6307
rect 21315 6273 21324 6307
rect 21272 6264 21324 6273
rect 22376 6264 22428 6316
rect 22560 6264 22612 6316
rect 22652 6307 22704 6316
rect 22652 6273 22661 6307
rect 22661 6273 22695 6307
rect 22695 6273 22704 6307
rect 22652 6264 22704 6273
rect 22744 6264 22796 6316
rect 22928 6307 22980 6316
rect 22928 6273 22937 6307
rect 22937 6273 22971 6307
rect 22971 6273 22980 6307
rect 22928 6264 22980 6273
rect 24124 6332 24176 6384
rect 21916 6196 21968 6248
rect 16580 6060 16632 6112
rect 19708 6103 19760 6112
rect 19708 6069 19717 6103
rect 19717 6069 19751 6103
rect 19751 6069 19760 6103
rect 19708 6060 19760 6069
rect 19800 6060 19852 6112
rect 19984 6103 20036 6112
rect 19984 6069 19993 6103
rect 19993 6069 20027 6103
rect 20027 6069 20036 6103
rect 19984 6060 20036 6069
rect 22008 6060 22060 6112
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 22376 6060 22428 6112
rect 4101 5958 4153 6010
rect 4165 5958 4217 6010
rect 4229 5958 4281 6010
rect 4293 5958 4345 6010
rect 4357 5958 4409 6010
rect 10403 5958 10455 6010
rect 10467 5958 10519 6010
rect 10531 5958 10583 6010
rect 10595 5958 10647 6010
rect 10659 5958 10711 6010
rect 16705 5958 16757 6010
rect 16769 5958 16821 6010
rect 16833 5958 16885 6010
rect 16897 5958 16949 6010
rect 16961 5958 17013 6010
rect 23007 5958 23059 6010
rect 23071 5958 23123 6010
rect 23135 5958 23187 6010
rect 23199 5958 23251 6010
rect 23263 5958 23315 6010
rect 3792 5856 3844 5908
rect 8116 5856 8168 5908
rect 6184 5788 6236 5840
rect 7196 5788 7248 5840
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 6000 5652 6052 5704
rect 6828 5652 6880 5704
rect 7564 5831 7616 5840
rect 7564 5797 7573 5831
rect 7573 5797 7607 5831
rect 7607 5797 7616 5831
rect 7564 5788 7616 5797
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 8576 5831 8628 5840
rect 8576 5797 8585 5831
rect 8585 5797 8619 5831
rect 8619 5797 8628 5831
rect 8576 5788 8628 5797
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 6092 5584 6144 5636
rect 9588 5788 9640 5840
rect 8852 5720 8904 5772
rect 9956 5856 10008 5908
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 11060 5856 11112 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 15568 5856 15620 5908
rect 17132 5856 17184 5908
rect 18604 5856 18656 5908
rect 20628 5856 20680 5908
rect 10784 5831 10836 5840
rect 10784 5797 10793 5831
rect 10793 5797 10827 5831
rect 10827 5797 10836 5831
rect 10784 5788 10836 5797
rect 11336 5831 11388 5840
rect 11336 5797 11345 5831
rect 11345 5797 11379 5831
rect 11379 5797 11388 5831
rect 11336 5788 11388 5797
rect 14096 5788 14148 5840
rect 12808 5720 12860 5772
rect 9772 5652 9824 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 8760 5584 8812 5636
rect 10784 5652 10836 5704
rect 12900 5652 12952 5704
rect 19524 5788 19576 5840
rect 21640 5856 21692 5908
rect 22928 5856 22980 5908
rect 15292 5652 15344 5704
rect 15384 5652 15436 5704
rect 15844 5720 15896 5772
rect 17776 5720 17828 5772
rect 21916 5720 21968 5772
rect 22560 5720 22612 5772
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 17960 5695 18012 5704
rect 17960 5661 17969 5695
rect 17969 5661 18003 5695
rect 18003 5661 18012 5695
rect 17960 5652 18012 5661
rect 20260 5652 20312 5704
rect 7656 5516 7708 5568
rect 8300 5516 8352 5568
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 11520 5516 11572 5568
rect 13176 5584 13228 5636
rect 17224 5584 17276 5636
rect 11980 5516 12032 5568
rect 14740 5559 14792 5568
rect 14740 5525 14765 5559
rect 14765 5525 14792 5559
rect 14740 5516 14792 5525
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 16396 5516 16448 5568
rect 16672 5516 16724 5568
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 22284 5652 22336 5704
rect 22744 5695 22796 5704
rect 22744 5661 22753 5695
rect 22753 5661 22787 5695
rect 22787 5661 22796 5695
rect 22744 5652 22796 5661
rect 20812 5584 20864 5636
rect 21732 5584 21784 5636
rect 22008 5584 22060 5636
rect 23572 5584 23624 5636
rect 22376 5516 22428 5568
rect 4761 5414 4813 5466
rect 4825 5414 4877 5466
rect 4889 5414 4941 5466
rect 4953 5414 5005 5466
rect 5017 5414 5069 5466
rect 11063 5414 11115 5466
rect 11127 5414 11179 5466
rect 11191 5414 11243 5466
rect 11255 5414 11307 5466
rect 11319 5414 11371 5466
rect 17365 5414 17417 5466
rect 17429 5414 17481 5466
rect 17493 5414 17545 5466
rect 17557 5414 17609 5466
rect 17621 5414 17673 5466
rect 23667 5414 23719 5466
rect 23731 5414 23783 5466
rect 23795 5414 23847 5466
rect 23859 5414 23911 5466
rect 23923 5414 23975 5466
rect 5724 5312 5776 5364
rect 7196 5355 7248 5364
rect 7196 5321 7221 5355
rect 7221 5321 7248 5355
rect 7196 5312 7248 5321
rect 6736 5244 6788 5296
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7840 5312 7892 5364
rect 11612 5312 11664 5364
rect 15200 5312 15252 5364
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 16488 5312 16540 5364
rect 15108 5244 15160 5296
rect 7564 5176 7616 5228
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 10324 5176 10376 5228
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 14924 5176 14976 5228
rect 17224 5312 17276 5364
rect 20260 5355 20312 5364
rect 20260 5321 20290 5355
rect 20290 5321 20312 5355
rect 20260 5312 20312 5321
rect 20996 5312 21048 5364
rect 17132 5244 17184 5296
rect 9496 5108 9548 5160
rect 10784 5108 10836 5160
rect 11060 5108 11112 5160
rect 14372 5108 14424 5160
rect 7932 5040 7984 5092
rect 7012 4972 7064 5024
rect 7564 4972 7616 5024
rect 10968 4972 11020 5024
rect 11152 4972 11204 5024
rect 11612 4972 11664 5024
rect 14188 4972 14240 5024
rect 14740 4972 14792 5024
rect 14924 4972 14976 5024
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 15936 5151 15988 5160
rect 15936 5117 15945 5151
rect 15945 5117 15979 5151
rect 15979 5117 15988 5151
rect 15936 5108 15988 5117
rect 16580 5108 16632 5160
rect 18052 5244 18104 5296
rect 19432 5244 19484 5296
rect 19524 5287 19576 5296
rect 19524 5253 19549 5287
rect 19549 5253 19576 5287
rect 19524 5244 19576 5253
rect 19984 5244 20036 5296
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 22008 5176 22060 5228
rect 22744 5312 22796 5364
rect 20444 5108 20496 5160
rect 22560 5176 22612 5228
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 16212 5040 16264 5092
rect 17040 5040 17092 5092
rect 16580 4972 16632 5024
rect 16672 4972 16724 5024
rect 17224 4972 17276 5024
rect 17960 5015 18012 5024
rect 17960 4981 17969 5015
rect 17969 4981 18003 5015
rect 18003 4981 18012 5015
rect 17960 4972 18012 4981
rect 19616 4972 19668 5024
rect 20076 4972 20128 5024
rect 22652 5083 22704 5092
rect 22652 5049 22661 5083
rect 22661 5049 22695 5083
rect 22695 5049 22704 5083
rect 22652 5040 22704 5049
rect 20812 4972 20864 5024
rect 4101 4870 4153 4922
rect 4165 4870 4217 4922
rect 4229 4870 4281 4922
rect 4293 4870 4345 4922
rect 4357 4870 4409 4922
rect 10403 4870 10455 4922
rect 10467 4870 10519 4922
rect 10531 4870 10583 4922
rect 10595 4870 10647 4922
rect 10659 4870 10711 4922
rect 16705 4870 16757 4922
rect 16769 4870 16821 4922
rect 16833 4870 16885 4922
rect 16897 4870 16949 4922
rect 16961 4870 17013 4922
rect 23007 4870 23059 4922
rect 23071 4870 23123 4922
rect 23135 4870 23187 4922
rect 23199 4870 23251 4922
rect 23263 4870 23315 4922
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 7840 4768 7892 4820
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 11060 4768 11112 4820
rect 5540 4564 5592 4616
rect 5724 4564 5776 4616
rect 6092 4564 6144 4616
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 7932 4564 7984 4616
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 11520 4700 11572 4752
rect 11704 4700 11756 4752
rect 14556 4700 14608 4752
rect 19432 4700 19484 4752
rect 20168 4743 20220 4752
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 11888 4632 11940 4684
rect 4620 4428 4672 4480
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 10048 4496 10100 4548
rect 6552 4471 6604 4480
rect 6552 4437 6561 4471
rect 6561 4437 6595 4471
rect 6595 4437 6604 4471
rect 6552 4428 6604 4437
rect 7656 4428 7708 4480
rect 7748 4471 7800 4480
rect 7748 4437 7757 4471
rect 7757 4437 7791 4471
rect 7791 4437 7800 4471
rect 7748 4428 7800 4437
rect 8392 4428 8444 4480
rect 10968 4428 11020 4480
rect 12624 4564 12676 4616
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 15016 4632 15068 4684
rect 20168 4709 20177 4743
rect 20177 4709 20211 4743
rect 20211 4709 20220 4743
rect 20168 4700 20220 4709
rect 19616 4675 19668 4684
rect 19616 4641 19625 4675
rect 19625 4641 19659 4675
rect 19659 4641 19668 4675
rect 19616 4632 19668 4641
rect 13912 4564 13964 4616
rect 14464 4607 14516 4616
rect 14464 4573 14467 4607
rect 14467 4573 14501 4607
rect 14501 4573 14516 4607
rect 14464 4564 14516 4573
rect 15292 4564 15344 4616
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 13636 4496 13688 4548
rect 14004 4496 14056 4548
rect 14740 4539 14792 4548
rect 14740 4505 14749 4539
rect 14749 4505 14783 4539
rect 14783 4505 14792 4539
rect 14740 4496 14792 4505
rect 14832 4496 14884 4548
rect 15936 4496 15988 4548
rect 17408 4564 17460 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20260 4675 20312 4684
rect 20260 4641 20269 4675
rect 20269 4641 20303 4675
rect 20303 4641 20312 4675
rect 20260 4632 20312 4641
rect 20444 4632 20496 4684
rect 20812 4675 20864 4684
rect 20812 4641 20821 4675
rect 20821 4641 20855 4675
rect 20855 4641 20864 4675
rect 20812 4632 20864 4641
rect 19984 4496 20036 4548
rect 14924 4428 14976 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 16856 4428 16908 4480
rect 19248 4471 19300 4480
rect 19248 4437 19257 4471
rect 19257 4437 19291 4471
rect 19291 4437 19300 4471
rect 19248 4428 19300 4437
rect 20260 4428 20312 4480
rect 21732 4675 21784 4684
rect 21732 4641 21741 4675
rect 21741 4641 21775 4675
rect 21775 4641 21784 4675
rect 21732 4632 21784 4641
rect 20996 4428 21048 4480
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 22008 4496 22060 4548
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 22376 4428 22428 4480
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 4761 4326 4813 4378
rect 4825 4326 4877 4378
rect 4889 4326 4941 4378
rect 4953 4326 5005 4378
rect 5017 4326 5069 4378
rect 11063 4326 11115 4378
rect 11127 4326 11179 4378
rect 11191 4326 11243 4378
rect 11255 4326 11307 4378
rect 11319 4326 11371 4378
rect 17365 4326 17417 4378
rect 17429 4326 17481 4378
rect 17493 4326 17545 4378
rect 17557 4326 17609 4378
rect 17621 4326 17673 4378
rect 23667 4326 23719 4378
rect 23731 4326 23783 4378
rect 23795 4326 23847 4378
rect 23859 4326 23911 4378
rect 23923 4326 23975 4378
rect 5540 4224 5592 4276
rect 4620 4199 4672 4208
rect 4620 4165 4654 4199
rect 4654 4165 4672 4199
rect 4620 4156 4672 4165
rect 7748 4224 7800 4276
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 6736 4156 6788 4208
rect 7104 4156 7156 4208
rect 5632 4088 5684 4140
rect 5448 4020 5500 4072
rect 6552 4020 6604 4072
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 7656 4199 7708 4208
rect 7656 4165 7665 4199
rect 7665 4165 7699 4199
rect 7699 4165 7708 4199
rect 7656 4156 7708 4165
rect 8208 4156 8260 4208
rect 7932 4088 7984 4140
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8392 4131 8444 4140
rect 8392 4097 8426 4131
rect 8426 4097 8444 4131
rect 8392 4088 8444 4097
rect 10048 4199 10100 4208
rect 10048 4165 10057 4199
rect 10057 4165 10091 4199
rect 10091 4165 10100 4199
rect 10048 4156 10100 4165
rect 9864 4088 9916 4140
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 13636 4224 13688 4276
rect 13728 4224 13780 4276
rect 14464 4224 14516 4276
rect 16488 4224 16540 4276
rect 17132 4224 17184 4276
rect 19984 4224 20036 4276
rect 20812 4224 20864 4276
rect 10784 4156 10836 4208
rect 11520 4199 11572 4208
rect 11520 4165 11529 4199
rect 11529 4165 11563 4199
rect 11563 4165 11572 4199
rect 11520 4156 11572 4165
rect 11612 4156 11664 4208
rect 14372 4156 14424 4208
rect 7104 4020 7156 4072
rect 9220 4020 9272 4072
rect 10968 4088 11020 4140
rect 11152 4088 11204 4140
rect 5540 3952 5592 4004
rect 5724 3952 5776 4004
rect 6368 3952 6420 4004
rect 6092 3884 6144 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 6644 3884 6696 3936
rect 6920 3952 6972 4004
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 12808 4088 12860 4140
rect 11152 3952 11204 4004
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 14280 4088 14332 4140
rect 17960 4156 18012 4208
rect 19340 4156 19392 4208
rect 14188 4063 14240 4072
rect 14188 4029 14197 4063
rect 14197 4029 14231 4063
rect 14231 4029 14240 4063
rect 14188 4020 14240 4029
rect 14832 4020 14884 4072
rect 15200 4088 15252 4140
rect 15844 4088 15896 4140
rect 15936 4088 15988 4140
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 16212 4063 16264 4072
rect 16212 4029 16221 4063
rect 16221 4029 16255 4063
rect 16255 4029 16264 4063
rect 16212 4020 16264 4029
rect 17132 4131 17184 4140
rect 17132 4097 17167 4131
rect 17167 4097 17184 4131
rect 17132 4088 17184 4097
rect 17776 4088 17828 4140
rect 20260 4088 20312 4140
rect 20536 4088 20588 4140
rect 22468 4156 22520 4208
rect 22928 4199 22980 4208
rect 22928 4165 22937 4199
rect 22937 4165 22971 4199
rect 22971 4165 22980 4199
rect 22928 4156 22980 4165
rect 21640 4088 21692 4140
rect 22376 4088 22428 4140
rect 22652 4131 22704 4140
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 19248 4020 19300 4072
rect 20076 4020 20128 4072
rect 19616 3952 19668 4004
rect 20996 4063 21048 4072
rect 20996 4029 21005 4063
rect 21005 4029 21039 4063
rect 21039 4029 21048 4063
rect 20996 4020 21048 4029
rect 22284 4063 22336 4072
rect 22284 4029 22293 4063
rect 22293 4029 22327 4063
rect 22327 4029 22336 4063
rect 22284 4020 22336 4029
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 8484 3884 8536 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 11060 3927 11112 3936
rect 11060 3893 11069 3927
rect 11069 3893 11103 3927
rect 11103 3893 11112 3927
rect 11060 3884 11112 3893
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 14372 3884 14424 3936
rect 14740 3884 14792 3936
rect 17040 3884 17092 3936
rect 22652 3884 22704 3936
rect 4101 3782 4153 3834
rect 4165 3782 4217 3834
rect 4229 3782 4281 3834
rect 4293 3782 4345 3834
rect 4357 3782 4409 3834
rect 10403 3782 10455 3834
rect 10467 3782 10519 3834
rect 10531 3782 10583 3834
rect 10595 3782 10647 3834
rect 10659 3782 10711 3834
rect 16705 3782 16757 3834
rect 16769 3782 16821 3834
rect 16833 3782 16885 3834
rect 16897 3782 16949 3834
rect 16961 3782 17013 3834
rect 23007 3782 23059 3834
rect 23071 3782 23123 3834
rect 23135 3782 23187 3834
rect 23199 3782 23251 3834
rect 23263 3782 23315 3834
rect 7840 3680 7892 3732
rect 9220 3680 9272 3732
rect 11980 3680 12032 3732
rect 12440 3680 12492 3732
rect 18236 3680 18288 3732
rect 20812 3680 20864 3732
rect 22376 3680 22428 3732
rect 6920 3612 6972 3664
rect 5540 3544 5592 3596
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 5448 3476 5500 3528
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 8116 3612 8168 3664
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 8668 3655 8720 3664
rect 8668 3621 8677 3655
rect 8677 3621 8711 3655
rect 8711 3621 8720 3655
rect 8668 3612 8720 3621
rect 14280 3612 14332 3664
rect 5632 3476 5684 3485
rect 7196 3476 7248 3528
rect 12900 3544 12952 3596
rect 14372 3587 14424 3596
rect 14372 3553 14381 3587
rect 14381 3553 14415 3587
rect 14415 3553 14424 3587
rect 14372 3544 14424 3553
rect 6000 3408 6052 3460
rect 7656 3408 7708 3460
rect 4620 3340 4672 3392
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 8208 3408 8260 3460
rect 9956 3476 10008 3528
rect 11060 3476 11112 3528
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 14096 3476 14148 3528
rect 14556 3476 14608 3528
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 8760 3408 8812 3460
rect 12992 3408 13044 3460
rect 13636 3408 13688 3460
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 17776 3612 17828 3664
rect 22652 3544 22704 3596
rect 24308 3680 24360 3732
rect 17132 3476 17184 3528
rect 18144 3476 18196 3528
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19340 3476 19392 3528
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 13084 3340 13136 3392
rect 14004 3340 14056 3392
rect 15752 3340 15804 3392
rect 16488 3340 16540 3392
rect 20444 3408 20496 3460
rect 21916 3408 21968 3460
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 19892 3340 19944 3392
rect 23572 3476 23624 3528
rect 4761 3238 4813 3290
rect 4825 3238 4877 3290
rect 4889 3238 4941 3290
rect 4953 3238 5005 3290
rect 5017 3238 5069 3290
rect 11063 3238 11115 3290
rect 11127 3238 11179 3290
rect 11191 3238 11243 3290
rect 11255 3238 11307 3290
rect 11319 3238 11371 3290
rect 17365 3238 17417 3290
rect 17429 3238 17481 3290
rect 17493 3238 17545 3290
rect 17557 3238 17609 3290
rect 17621 3238 17673 3290
rect 23667 3238 23719 3290
rect 23731 3238 23783 3290
rect 23795 3238 23847 3290
rect 23859 3238 23911 3290
rect 23923 3238 23975 3290
rect 5816 3136 5868 3188
rect 6736 3136 6788 3188
rect 8760 3136 8812 3188
rect 11612 3136 11664 3188
rect 15200 3136 15252 3188
rect 17868 3136 17920 3188
rect 20260 3179 20312 3188
rect 20260 3145 20269 3179
rect 20269 3145 20303 3179
rect 20303 3145 20312 3179
rect 20260 3136 20312 3145
rect 20444 3179 20496 3188
rect 20444 3145 20453 3179
rect 20453 3145 20487 3179
rect 20487 3145 20496 3179
rect 20444 3136 20496 3145
rect 21916 3136 21968 3188
rect 5632 3068 5684 3120
rect 6368 3111 6420 3120
rect 6368 3077 6377 3111
rect 6377 3077 6411 3111
rect 6411 3077 6420 3111
rect 6368 3068 6420 3077
rect 10048 3068 10100 3120
rect 13820 3068 13872 3120
rect 18144 3068 18196 3120
rect 18604 3068 18656 3120
rect 4620 2932 4672 2984
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 12900 2932 12952 2984
rect 17040 2975 17092 2984
rect 17040 2941 17049 2975
rect 17049 2941 17083 2975
rect 17083 2941 17092 2975
rect 17040 2932 17092 2941
rect 19892 3000 19944 3052
rect 20812 3068 20864 3120
rect 17776 2932 17828 2984
rect 18880 2932 18932 2984
rect 21180 3000 21232 3052
rect 20168 2932 20220 2984
rect 6644 2907 6696 2916
rect 6644 2873 6653 2907
rect 6653 2873 6687 2907
rect 6687 2873 6696 2907
rect 6644 2864 6696 2873
rect 19432 2864 19484 2916
rect 4101 2694 4153 2746
rect 4165 2694 4217 2746
rect 4229 2694 4281 2746
rect 4293 2694 4345 2746
rect 4357 2694 4409 2746
rect 10403 2694 10455 2746
rect 10467 2694 10519 2746
rect 10531 2694 10583 2746
rect 10595 2694 10647 2746
rect 10659 2694 10711 2746
rect 16705 2694 16757 2746
rect 16769 2694 16821 2746
rect 16833 2694 16885 2746
rect 16897 2694 16949 2746
rect 16961 2694 17013 2746
rect 23007 2694 23059 2746
rect 23071 2694 23123 2746
rect 23135 2694 23187 2746
rect 23199 2694 23251 2746
rect 23263 2694 23315 2746
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 9128 2592 9180 2644
rect 12072 2592 12124 2644
rect 13820 2635 13872 2644
rect 13820 2601 13829 2635
rect 13829 2601 13863 2635
rect 13863 2601 13872 2635
rect 13820 2592 13872 2601
rect 16304 2592 16356 2644
rect 23572 2592 23624 2644
rect 11428 2456 11480 2508
rect 3884 2388 3936 2440
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 7748 2388 7800 2440
rect 11612 2388 11664 2440
rect 12808 2388 12860 2440
rect 17132 2524 17184 2576
rect 14464 2456 14516 2508
rect 15476 2388 15528 2440
rect 24032 2388 24084 2440
rect 20 2320 72 2372
rect 13452 2320 13504 2372
rect 10876 2252 10928 2304
rect 19984 2252 20036 2304
rect 24768 2252 24820 2304
rect 4761 2150 4813 2202
rect 4825 2150 4877 2202
rect 4889 2150 4941 2202
rect 4953 2150 5005 2202
rect 5017 2150 5069 2202
rect 11063 2150 11115 2202
rect 11127 2150 11179 2202
rect 11191 2150 11243 2202
rect 11255 2150 11307 2202
rect 11319 2150 11371 2202
rect 17365 2150 17417 2202
rect 17429 2150 17481 2202
rect 17493 2150 17545 2202
rect 17557 2150 17609 2202
rect 17621 2150 17673 2202
rect 23667 2150 23719 2202
rect 23731 2150 23783 2202
rect 23795 2150 23847 2202
rect 23859 2150 23911 2202
rect 23923 2150 23975 2202
<< metal2 >>
rect 1398 29336 1454 29345
rect 1398 29271 1454 29280
rect 1412 26994 1440 29271
rect 3238 28825 3294 29625
rect 7102 28825 7158 29625
rect 11610 28825 11666 29625
rect 15474 28825 15530 29625
rect 19338 28825 19394 29625
rect 23202 28825 23258 29625
rect 27066 28825 27122 29625
rect 3252 27130 3280 28825
rect 4761 27228 5069 27237
rect 4761 27226 4767 27228
rect 4823 27226 4847 27228
rect 4903 27226 4927 27228
rect 4983 27226 5007 27228
rect 5063 27226 5069 27228
rect 4823 27174 4825 27226
rect 5005 27174 5007 27226
rect 4761 27172 4767 27174
rect 4823 27172 4847 27174
rect 4903 27172 4927 27174
rect 4983 27172 5007 27174
rect 5063 27172 5069 27174
rect 4761 27163 5069 27172
rect 7116 27130 7144 28825
rect 11063 27228 11371 27237
rect 11063 27226 11069 27228
rect 11125 27226 11149 27228
rect 11205 27226 11229 27228
rect 11285 27226 11309 27228
rect 11365 27226 11371 27228
rect 11125 27174 11127 27226
rect 11307 27174 11309 27226
rect 11063 27172 11069 27174
rect 11125 27172 11149 27174
rect 11205 27172 11229 27174
rect 11285 27172 11309 27174
rect 11365 27172 11371 27174
rect 11063 27163 11371 27172
rect 11624 27130 11652 28825
rect 3240 27124 3292 27130
rect 3240 27066 3292 27072
rect 7104 27124 7156 27130
rect 7104 27066 7156 27072
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 10784 27056 10836 27062
rect 10784 26998 10836 27004
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 2596 26784 2648 26790
rect 2596 26726 2648 26732
rect 2504 21616 2556 21622
rect 2504 21558 2556 21564
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 952 20942 980 21111
rect 940 20936 992 20942
rect 940 20878 992 20884
rect 1412 19378 1440 21422
rect 2148 21146 2176 21422
rect 2516 21146 2544 21558
rect 2136 21140 2188 21146
rect 2136 21082 2188 21088
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1596 20505 1624 20742
rect 1582 20496 1638 20505
rect 1582 20431 1638 20440
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19446 1716 19654
rect 1676 19440 1728 19446
rect 1676 19382 1728 19388
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 2332 18766 2360 20878
rect 2608 19825 2636 26726
rect 4101 26684 4409 26693
rect 4101 26682 4107 26684
rect 4163 26682 4187 26684
rect 4243 26682 4267 26684
rect 4323 26682 4347 26684
rect 4403 26682 4409 26684
rect 4163 26630 4165 26682
rect 4345 26630 4347 26682
rect 4101 26628 4107 26630
rect 4163 26628 4187 26630
rect 4243 26628 4267 26630
rect 4323 26628 4347 26630
rect 4403 26628 4409 26630
rect 4101 26619 4409 26628
rect 10403 26684 10711 26693
rect 10403 26682 10409 26684
rect 10465 26682 10489 26684
rect 10545 26682 10569 26684
rect 10625 26682 10649 26684
rect 10705 26682 10711 26684
rect 10465 26630 10467 26682
rect 10647 26630 10649 26682
rect 10403 26628 10409 26630
rect 10465 26628 10489 26630
rect 10545 26628 10569 26630
rect 10625 26628 10649 26630
rect 10705 26628 10711 26630
rect 10403 26619 10711 26628
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 6552 26376 6604 26382
rect 6552 26318 6604 26324
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 4761 26140 5069 26149
rect 4761 26138 4767 26140
rect 4823 26138 4847 26140
rect 4903 26138 4927 26140
rect 4983 26138 5007 26140
rect 5063 26138 5069 26140
rect 4823 26086 4825 26138
rect 5005 26086 5007 26138
rect 4761 26084 4767 26086
rect 4823 26084 4847 26086
rect 4903 26084 4927 26086
rect 4983 26084 5007 26086
rect 5063 26084 5069 26086
rect 4761 26075 5069 26084
rect 6564 25974 6592 26318
rect 7472 26308 7524 26314
rect 7472 26250 7524 26256
rect 6552 25968 6604 25974
rect 6552 25910 6604 25916
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 4101 25596 4409 25605
rect 4101 25594 4107 25596
rect 4163 25594 4187 25596
rect 4243 25594 4267 25596
rect 4323 25594 4347 25596
rect 4403 25594 4409 25596
rect 4163 25542 4165 25594
rect 4345 25542 4347 25594
rect 4101 25540 4107 25542
rect 4163 25540 4187 25542
rect 4243 25540 4267 25542
rect 4323 25540 4347 25542
rect 4403 25540 4409 25542
rect 4101 25531 4409 25540
rect 6564 25362 6592 25910
rect 6932 25498 6960 25910
rect 7484 25498 7512 26250
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 8312 25362 8340 26182
rect 8956 25974 8984 26318
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 8944 25968 8996 25974
rect 8864 25928 8944 25956
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 3238 25256 3294 25265
rect 3238 25191 3294 25200
rect 6000 25220 6052 25226
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2780 21140 2832 21146
rect 2780 21082 2832 21088
rect 2792 19854 2820 21082
rect 2884 21010 2912 21354
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 2884 20466 2912 20946
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2884 20058 2912 20198
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19848 2832 19854
rect 2594 19816 2650 19825
rect 2780 19790 2832 19796
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2594 19751 2650 19760
rect 2976 19514 3004 19790
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2792 18970 2820 19314
rect 3160 19310 3188 20402
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 940 16584 992 16590
rect 940 16526 992 16532
rect 952 16425 980 16526
rect 938 16416 994 16425
rect 938 16351 994 16360
rect 1412 15570 1440 17614
rect 1688 17610 1716 18022
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 2332 17202 2360 18702
rect 3252 18358 3280 25191
rect 6000 25162 6052 25168
rect 4761 25052 5069 25061
rect 4761 25050 4767 25052
rect 4823 25050 4847 25052
rect 4903 25050 4927 25052
rect 4983 25050 5007 25052
rect 5063 25050 5069 25052
rect 4823 24998 4825 25050
rect 5005 24998 5007 25050
rect 4761 24996 4767 24998
rect 4823 24996 4847 24998
rect 4903 24996 4927 24998
rect 4983 24996 5007 24998
rect 5063 24996 5069 24998
rect 4761 24987 5069 24996
rect 6012 24818 6040 25162
rect 6564 25158 6592 25298
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6736 25220 6788 25226
rect 6736 25162 6788 25168
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 6000 24812 6052 24818
rect 6000 24754 6052 24760
rect 4101 24508 4409 24517
rect 4101 24506 4107 24508
rect 4163 24506 4187 24508
rect 4243 24506 4267 24508
rect 4323 24506 4347 24508
rect 4403 24506 4409 24508
rect 4163 24454 4165 24506
rect 4345 24454 4347 24506
rect 4101 24452 4107 24454
rect 4163 24452 4187 24454
rect 4243 24452 4267 24454
rect 4323 24452 4347 24454
rect 4403 24452 4409 24454
rect 4101 24443 4409 24452
rect 6472 24410 6500 25094
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6564 24274 6592 25094
rect 6748 24818 6776 25162
rect 6840 24886 6868 25230
rect 8772 25226 8800 25774
rect 8760 25220 8812 25226
rect 8760 25162 8812 25168
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 6828 24880 6880 24886
rect 6828 24822 6880 24828
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6000 24200 6052 24206
rect 6000 24142 6052 24148
rect 4761 23964 5069 23973
rect 4761 23962 4767 23964
rect 4823 23962 4847 23964
rect 4903 23962 4927 23964
rect 4983 23962 5007 23964
rect 5063 23962 5069 23964
rect 4823 23910 4825 23962
rect 5005 23910 5007 23962
rect 4761 23908 4767 23910
rect 4823 23908 4847 23910
rect 4903 23908 4927 23910
rect 4983 23908 5007 23910
rect 5063 23908 5069 23910
rect 4761 23899 5069 23908
rect 6012 23798 6040 24142
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6564 23866 6592 24074
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 3700 23792 3752 23798
rect 5172 23792 5224 23798
rect 3700 23734 3752 23740
rect 5170 23760 5172 23769
rect 6000 23792 6052 23798
rect 5224 23760 5226 23769
rect 3712 23526 3740 23734
rect 6000 23734 6052 23740
rect 5170 23695 5226 23704
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6472 23633 6500 23666
rect 6840 23633 6868 24822
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 7472 24676 7524 24682
rect 7472 24618 7524 24624
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7300 23730 7328 24550
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 6458 23624 6514 23633
rect 5540 23588 5592 23594
rect 6458 23559 6514 23568
rect 6826 23624 6882 23633
rect 7484 23594 7512 24618
rect 7576 23662 7604 24754
rect 7668 24070 7696 24754
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7668 23594 7696 24006
rect 7760 23866 7788 24006
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7852 23798 7880 24754
rect 8036 24682 8064 24754
rect 8024 24676 8076 24682
rect 8024 24618 8076 24624
rect 8036 24410 8064 24618
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 8128 24188 8156 24890
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8220 24342 8248 24550
rect 8208 24336 8260 24342
rect 8208 24278 8260 24284
rect 8208 24200 8260 24206
rect 8128 24160 8208 24188
rect 8208 24142 8260 24148
rect 8312 24070 8340 24686
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8496 24138 8524 24550
rect 8588 24410 8800 24426
rect 8576 24404 8800 24410
rect 8628 24398 8800 24404
rect 8576 24346 8628 24352
rect 8392 24132 8444 24138
rect 8392 24074 8444 24080
rect 8484 24132 8536 24138
rect 8484 24074 8536 24080
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 7840 23792 7892 23798
rect 7840 23734 7892 23740
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 6826 23559 6882 23568
rect 7472 23588 7524 23594
rect 5540 23530 5592 23536
rect 3700 23520 3752 23526
rect 5552 23497 5580 23530
rect 5632 23520 5684 23526
rect 3700 23462 3752 23468
rect 5538 23488 5594 23497
rect 3608 23112 3660 23118
rect 3608 23054 3660 23060
rect 3620 21690 3648 23054
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3516 21616 3568 21622
rect 3516 21558 3568 21564
rect 3528 21146 3556 21558
rect 3620 21554 3648 21626
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3620 21350 3648 21490
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3332 21004 3384 21010
rect 3332 20946 3384 20952
rect 3344 19854 3372 20946
rect 3436 20602 3464 21082
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3436 19854 3464 19994
rect 3528 19922 3556 20334
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3436 19174 3464 19790
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3620 18222 3648 19110
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3068 17678 3096 18158
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2424 17338 2452 17546
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2148 16794 2176 17138
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2332 16250 2360 17138
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 2228 15904 2280 15910
rect 2228 15846 2280 15852
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 15162 1440 15506
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1412 15026 1440 15098
rect 1688 15094 1716 15846
rect 2240 15570 2268 15846
rect 2332 15706 2360 16050
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 1676 15088 1728 15094
rect 1676 15030 1728 15036
rect 2792 15026 2820 15914
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15502 3004 15846
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 9110 1808 9522
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1768 9104 1820 9110
rect 1768 9046 1820 9052
rect 1872 9042 1900 9454
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1964 8634 1992 14282
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2148 12306 2176 12718
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11830 2084 12038
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 2148 10198 2176 12242
rect 2240 11626 2268 12786
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2424 10742 2452 11834
rect 2516 11626 2544 12106
rect 2700 11778 2728 12106
rect 2608 11762 2820 11778
rect 3068 11762 3096 12378
rect 2596 11756 2832 11762
rect 2648 11750 2780 11756
rect 2596 11698 2648 11704
rect 2780 11698 2832 11704
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2148 9586 2176 10134
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 9178 2360 9522
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2424 9058 2452 10678
rect 2608 10470 2636 11698
rect 3068 11354 3096 11698
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3252 11150 3280 11698
rect 3344 11286 3372 17614
rect 3620 17610 3648 18022
rect 3608 17604 3660 17610
rect 3608 17546 3660 17552
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12986 3556 13126
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3436 11762 3464 12378
rect 3528 12306 3556 12922
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2332 9030 2452 9058
rect 2332 8906 2360 9030
rect 2516 8906 2544 9318
rect 2608 9178 2636 10406
rect 2792 10062 2820 10406
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2884 9178 2912 10678
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 2332 8430 2360 8842
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2608 8294 2636 9114
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2700 8362 2728 8978
rect 3436 8974 3464 9318
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2596 8288 2648 8294
rect 1398 8256 1454 8265
rect 2596 8230 2648 8236
rect 1398 8191 1454 8200
rect 2608 8090 2636 8230
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2700 7954 2728 8298
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 3252 7818 3280 8434
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3620 7410 3648 7686
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3712 4185 3740 23462
rect 5632 23462 5684 23468
rect 4101 23420 4409 23429
rect 5538 23423 5594 23432
rect 4101 23418 4107 23420
rect 4163 23418 4187 23420
rect 4243 23418 4267 23420
rect 4323 23418 4347 23420
rect 4403 23418 4409 23420
rect 4163 23366 4165 23418
rect 4345 23366 4347 23418
rect 4101 23364 4107 23366
rect 4163 23364 4187 23366
rect 4243 23364 4267 23366
rect 4323 23364 4347 23366
rect 4403 23364 4409 23366
rect 4101 23355 4409 23364
rect 5644 23322 5672 23462
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 4068 23044 4120 23050
rect 4068 22986 4120 22992
rect 4080 22778 4108 22986
rect 4761 22876 5069 22885
rect 4761 22874 4767 22876
rect 4823 22874 4847 22876
rect 4903 22874 4927 22876
rect 4983 22874 5007 22876
rect 5063 22874 5069 22876
rect 4823 22822 4825 22874
rect 5005 22822 5007 22874
rect 4761 22820 4767 22822
rect 4823 22820 4847 22822
rect 4903 22820 4927 22822
rect 4983 22820 5007 22822
rect 5063 22820 5069 22822
rect 4761 22811 5069 22820
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 6012 22710 6040 23054
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6288 22778 6316 22918
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6000 22704 6052 22710
rect 6000 22646 6052 22652
rect 6472 22642 6500 23559
rect 7472 23530 7524 23536
rect 7656 23588 7708 23594
rect 7656 23530 7708 23536
rect 8220 23526 8248 23734
rect 8404 23594 8432 24074
rect 8496 23730 8524 24074
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8772 23594 8800 24398
rect 8864 24342 8892 25928
rect 8944 25910 8996 25916
rect 9128 25900 9180 25906
rect 9048 25860 9128 25888
rect 9048 25498 9076 25860
rect 9128 25842 9180 25848
rect 9232 25838 9260 26250
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9416 25702 9444 26250
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 9600 25974 9628 26182
rect 9588 25968 9640 25974
rect 9588 25910 9640 25916
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 9048 24818 9076 25434
rect 9128 25288 9180 25294
rect 9126 25256 9128 25265
rect 9180 25256 9182 25265
rect 9126 25191 9182 25200
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8852 24336 8904 24342
rect 8852 24278 8904 24284
rect 8864 24206 8892 24278
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8864 23866 8892 24142
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 8956 23730 8984 24550
rect 9048 24274 9076 24754
rect 9232 24614 9260 25638
rect 9416 25378 9444 25638
rect 9324 25350 9444 25378
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9036 24268 9088 24274
rect 9036 24210 9088 24216
rect 9232 23730 9260 24550
rect 9324 24410 9352 25350
rect 9600 25294 9628 25774
rect 9692 25294 9720 26454
rect 9864 26444 9916 26450
rect 9864 26386 9916 26392
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 25362 9812 26182
rect 9876 25430 9904 26386
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9968 25498 9996 26318
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10612 25906 10640 26250
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10232 25696 10284 25702
rect 10232 25638 10284 25644
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9864 25424 9916 25430
rect 9864 25366 9916 25372
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9404 25220 9456 25226
rect 9404 25162 9456 25168
rect 9416 24954 9444 25162
rect 9404 24948 9456 24954
rect 9404 24890 9456 24896
rect 9508 24732 9536 25230
rect 9968 25226 9996 25434
rect 10244 25430 10272 25638
rect 10403 25596 10711 25605
rect 10403 25594 10409 25596
rect 10465 25594 10489 25596
rect 10545 25594 10569 25596
rect 10625 25594 10649 25596
rect 10705 25594 10711 25596
rect 10465 25542 10467 25594
rect 10647 25542 10649 25594
rect 10403 25540 10409 25542
rect 10465 25540 10489 25542
rect 10545 25540 10569 25542
rect 10625 25540 10649 25542
rect 10705 25540 10711 25542
rect 10403 25531 10711 25540
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10232 25288 10284 25294
rect 10138 25256 10194 25265
rect 9956 25220 10008 25226
rect 10232 25230 10284 25236
rect 10138 25191 10194 25200
rect 9956 25162 10008 25168
rect 10152 24818 10180 25191
rect 10244 25158 10272 25230
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 9680 24744 9732 24750
rect 9508 24704 9680 24732
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9324 24206 9352 24346
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9404 24200 9456 24206
rect 9404 24142 9456 24148
rect 9310 23896 9366 23905
rect 9416 23866 9444 24142
rect 9508 24070 9536 24704
rect 9680 24686 9732 24692
rect 9680 24608 9732 24614
rect 9600 24568 9680 24596
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9310 23831 9366 23840
rect 9404 23860 9456 23866
rect 9324 23798 9352 23831
rect 9404 23802 9456 23808
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9508 23730 9536 24006
rect 9600 23798 9628 24568
rect 9680 24550 9732 24556
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9588 23792 9640 23798
rect 9588 23734 9640 23740
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 8392 23588 8444 23594
rect 8392 23530 8444 23536
rect 8760 23588 8812 23594
rect 8760 23530 8812 23536
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 9048 23322 9076 23598
rect 9128 23588 9180 23594
rect 9128 23530 9180 23536
rect 9496 23588 9548 23594
rect 9496 23530 9548 23536
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9140 23186 9168 23530
rect 9508 23497 9536 23530
rect 9494 23488 9550 23497
rect 9494 23423 9550 23432
rect 9128 23180 9180 23186
rect 9128 23122 9180 23128
rect 9600 23118 9628 23598
rect 9876 23322 9904 24142
rect 9956 24064 10008 24070
rect 9954 24032 9956 24041
rect 10008 24032 10010 24041
rect 9954 23967 10010 23976
rect 9968 23730 9996 23967
rect 10046 23896 10102 23905
rect 10046 23831 10102 23840
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 10060 23526 10088 23831
rect 10152 23798 10180 24754
rect 10244 24274 10272 25094
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 10152 23594 10180 23734
rect 10336 23730 10364 24618
rect 10403 24508 10711 24517
rect 10403 24506 10409 24508
rect 10465 24506 10489 24508
rect 10545 24506 10569 24508
rect 10625 24506 10649 24508
rect 10705 24506 10711 24508
rect 10465 24454 10467 24506
rect 10647 24454 10649 24506
rect 10403 24452 10409 24454
rect 10465 24452 10489 24454
rect 10545 24452 10569 24454
rect 10625 24452 10649 24454
rect 10705 24452 10711 24454
rect 10403 24443 10711 24452
rect 10690 24032 10746 24041
rect 10690 23967 10746 23976
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10704 23662 10732 23967
rect 10796 23746 10824 26998
rect 15488 26994 15516 28825
rect 17365 27228 17673 27237
rect 17365 27226 17371 27228
rect 17427 27226 17451 27228
rect 17507 27226 17531 27228
rect 17587 27226 17611 27228
rect 17667 27226 17673 27228
rect 17427 27174 17429 27226
rect 17609 27174 17611 27226
rect 17365 27172 17371 27174
rect 17427 27172 17451 27174
rect 17507 27172 17531 27174
rect 17587 27172 17611 27174
rect 17667 27172 17673 27174
rect 17365 27163 17673 27172
rect 19352 27130 19380 28825
rect 23216 27554 23244 28825
rect 23216 27526 23520 27554
rect 23492 27130 23520 27526
rect 23667 27228 23975 27237
rect 23667 27226 23673 27228
rect 23729 27226 23753 27228
rect 23809 27226 23833 27228
rect 23889 27226 23913 27228
rect 23969 27226 23975 27228
rect 23729 27174 23731 27226
rect 23911 27174 23913 27226
rect 23667 27172 23673 27174
rect 23729 27172 23753 27174
rect 23809 27172 23833 27174
rect 23889 27172 23913 27174
rect 23969 27172 23975 27174
rect 23667 27163 23975 27172
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 10876 26240 10928 26246
rect 10876 26182 10928 26188
rect 10888 25362 10916 26182
rect 11063 26140 11371 26149
rect 11063 26138 11069 26140
rect 11125 26138 11149 26140
rect 11205 26138 11229 26140
rect 11285 26138 11309 26140
rect 11365 26138 11371 26140
rect 11125 26086 11127 26138
rect 11307 26086 11309 26138
rect 11063 26084 11069 26086
rect 11125 26084 11149 26086
rect 11205 26084 11229 26086
rect 11285 26084 11309 26086
rect 11365 26084 11371 26086
rect 11063 26075 11371 26084
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 11063 25052 11371 25061
rect 11063 25050 11069 25052
rect 11125 25050 11149 25052
rect 11205 25050 11229 25052
rect 11285 25050 11309 25052
rect 11365 25050 11371 25052
rect 11125 24998 11127 25050
rect 11307 24998 11309 25050
rect 11063 24996 11069 24998
rect 11125 24996 11149 24998
rect 11205 24996 11229 24998
rect 11285 24996 11309 24998
rect 11365 24996 11371 24998
rect 11063 24987 11371 24996
rect 11063 23964 11371 23973
rect 11063 23962 11069 23964
rect 11125 23962 11149 23964
rect 11205 23962 11229 23964
rect 11285 23962 11309 23964
rect 11365 23962 11371 23964
rect 11125 23910 11127 23962
rect 11307 23910 11309 23962
rect 11063 23908 11069 23910
rect 11125 23908 11149 23910
rect 11205 23908 11229 23910
rect 11285 23908 11309 23910
rect 11365 23908 11371 23910
rect 11063 23899 11371 23908
rect 10796 23718 10916 23746
rect 10692 23656 10744 23662
rect 10692 23598 10744 23604
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10140 23588 10192 23594
rect 10140 23530 10192 23536
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 10048 23520 10100 23526
rect 10152 23497 10180 23530
rect 10704 23526 10732 23598
rect 10692 23520 10744 23526
rect 10048 23462 10100 23468
rect 10138 23488 10194 23497
rect 9968 23361 9996 23462
rect 9954 23352 10010 23361
rect 9772 23316 9824 23322
rect 9772 23258 9824 23264
rect 9864 23316 9916 23322
rect 9954 23287 10010 23296
rect 9864 23258 9916 23264
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9784 22710 9812 23258
rect 9956 23248 10008 23254
rect 9956 23190 10008 23196
rect 9968 22778 9996 23190
rect 10060 23118 10088 23462
rect 10692 23462 10744 23468
rect 10138 23423 10194 23432
rect 10403 23420 10711 23429
rect 10403 23418 10409 23420
rect 10465 23418 10489 23420
rect 10545 23418 10569 23420
rect 10625 23418 10649 23420
rect 10705 23418 10711 23420
rect 10465 23366 10467 23418
rect 10647 23366 10649 23418
rect 10403 23364 10409 23366
rect 10465 23364 10489 23366
rect 10545 23364 10569 23366
rect 10625 23364 10649 23366
rect 10705 23364 10711 23366
rect 10403 23355 10711 23364
rect 10796 23225 10824 23598
rect 10782 23216 10838 23225
rect 10782 23151 10838 23160
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10796 22778 10824 23151
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 9220 22704 9272 22710
rect 9220 22646 9272 22652
rect 9404 22704 9456 22710
rect 9404 22646 9456 22652
rect 9772 22704 9824 22710
rect 10888 22658 10916 23718
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11072 23633 11100 23666
rect 11058 23624 11114 23633
rect 11058 23559 11114 23568
rect 11063 22876 11371 22885
rect 11063 22874 11069 22876
rect 11125 22874 11149 22876
rect 11205 22874 11229 22876
rect 11285 22874 11309 22876
rect 11365 22874 11371 22876
rect 11125 22822 11127 22874
rect 11307 22822 11309 22874
rect 11063 22820 11069 22822
rect 11125 22820 11149 22822
rect 11205 22820 11229 22822
rect 11285 22820 11309 22822
rect 11365 22820 11371 22822
rect 11063 22811 11371 22820
rect 9772 22646 9824 22652
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 4101 22332 4409 22341
rect 4101 22330 4107 22332
rect 4163 22330 4187 22332
rect 4243 22330 4267 22332
rect 4323 22330 4347 22332
rect 4403 22330 4409 22332
rect 4163 22278 4165 22330
rect 4345 22278 4347 22330
rect 4101 22276 4107 22278
rect 4163 22276 4187 22278
rect 4243 22276 4267 22278
rect 4323 22276 4347 22278
rect 4403 22276 4409 22278
rect 4101 22267 4409 22276
rect 4160 22024 4212 22030
rect 4158 21992 4160 22001
rect 4908 22001 4936 22578
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 5724 22024 5776 22030
rect 4212 21992 4214 22001
rect 4158 21927 4214 21936
rect 4894 21992 4950 22001
rect 5724 21966 5776 21972
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 4894 21927 4950 21936
rect 3792 21888 3844 21894
rect 3792 21830 3844 21836
rect 3804 18426 3832 21830
rect 4761 21788 5069 21797
rect 4761 21786 4767 21788
rect 4823 21786 4847 21788
rect 4903 21786 4927 21788
rect 4983 21786 5007 21788
rect 5063 21786 5069 21788
rect 4823 21734 4825 21786
rect 5005 21734 5007 21786
rect 4761 21732 4767 21734
rect 4823 21732 4847 21734
rect 4903 21732 4927 21734
rect 4983 21732 5007 21734
rect 5063 21732 5069 21734
rect 4761 21723 5069 21732
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5552 21434 5580 21626
rect 5632 21480 5684 21486
rect 5552 21428 5632 21434
rect 5552 21422 5684 21428
rect 3896 21146 3924 21422
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3884 21140 3936 21146
rect 3884 21082 3936 21088
rect 3988 20942 4016 21286
rect 4101 21244 4409 21253
rect 4101 21242 4107 21244
rect 4163 21242 4187 21244
rect 4243 21242 4267 21244
rect 4323 21242 4347 21244
rect 4403 21242 4409 21244
rect 4163 21190 4165 21242
rect 4345 21190 4347 21242
rect 4101 21188 4107 21190
rect 4163 21188 4187 21190
rect 4243 21188 4267 21190
rect 4323 21188 4347 21190
rect 4403 21188 4409 21190
rect 4101 21179 4409 21188
rect 4344 21140 4396 21146
rect 4344 21082 4396 21088
rect 4356 20942 4384 21082
rect 5184 21078 5212 21422
rect 5552 21406 5672 21422
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4356 20466 4384 20878
rect 4344 20460 4396 20466
rect 4344 20402 4396 20408
rect 4448 20262 4476 20878
rect 4761 20700 5069 20709
rect 4761 20698 4767 20700
rect 4823 20698 4847 20700
rect 4903 20698 4927 20700
rect 4983 20698 5007 20700
rect 5063 20698 5069 20700
rect 4823 20646 4825 20698
rect 5005 20646 5007 20698
rect 4761 20644 4767 20646
rect 4823 20644 4847 20646
rect 4903 20644 4927 20646
rect 4983 20644 5007 20646
rect 5063 20644 5069 20646
rect 4761 20635 5069 20644
rect 5184 20534 5212 21014
rect 5276 20942 5304 21082
rect 5552 21010 5580 21406
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4101 20156 4409 20165
rect 4101 20154 4107 20156
rect 4163 20154 4187 20156
rect 4243 20154 4267 20156
rect 4323 20154 4347 20156
rect 4403 20154 4409 20156
rect 4163 20102 4165 20154
rect 4345 20102 4347 20154
rect 4101 20100 4107 20102
rect 4163 20100 4187 20102
rect 4243 20100 4267 20102
rect 4323 20100 4347 20102
rect 4403 20100 4409 20102
rect 4101 20091 4409 20100
rect 4448 20058 4476 20198
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 4448 19802 4476 19994
rect 4356 19774 4476 19802
rect 4356 19310 4384 19774
rect 4540 19718 4568 20198
rect 4724 19854 4752 20198
rect 4816 20058 4844 20402
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 5184 19922 5212 20470
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 4712 19848 4764 19854
rect 4632 19808 4712 19836
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 4448 19514 4476 19654
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4436 19236 4488 19242
rect 4436 19178 4488 19184
rect 4101 19068 4409 19077
rect 4101 19066 4107 19068
rect 4163 19066 4187 19068
rect 4243 19066 4267 19068
rect 4323 19066 4347 19068
rect 4403 19066 4409 19068
rect 4163 19014 4165 19066
rect 4345 19014 4347 19066
rect 4101 19012 4107 19014
rect 4163 19012 4187 19014
rect 4243 19012 4267 19014
rect 4323 19012 4347 19014
rect 4403 19012 4409 19014
rect 4101 19003 4409 19012
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3804 16250 3832 18362
rect 4448 18222 4476 19178
rect 4540 18272 4568 19654
rect 4632 19446 4660 19808
rect 4712 19790 4764 19796
rect 4761 19612 5069 19621
rect 4761 19610 4767 19612
rect 4823 19610 4847 19612
rect 4903 19610 4927 19612
rect 4983 19610 5007 19612
rect 5063 19610 5069 19612
rect 4823 19558 4825 19610
rect 5005 19558 5007 19610
rect 4761 19556 4767 19558
rect 4823 19556 4847 19558
rect 4903 19556 4927 19558
rect 4983 19556 5007 19558
rect 5063 19556 5069 19558
rect 4761 19547 5069 19556
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4620 19440 4672 19446
rect 4816 19417 4844 19450
rect 4620 19382 4672 19388
rect 4802 19408 4858 19417
rect 4632 19174 4660 19382
rect 5184 19378 5212 19858
rect 4802 19343 4858 19352
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 5276 18834 5304 20538
rect 5552 20466 5580 20742
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 20058 5396 20198
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5460 19922 5488 20334
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 4761 18524 5069 18533
rect 4761 18522 4767 18524
rect 4823 18522 4847 18524
rect 4903 18522 4927 18524
rect 4983 18522 5007 18524
rect 5063 18522 5069 18524
rect 4823 18470 4825 18522
rect 5005 18470 5007 18522
rect 4761 18468 4767 18470
rect 4823 18468 4847 18470
rect 4903 18468 4927 18470
rect 4983 18468 5007 18470
rect 5063 18468 5069 18470
rect 4761 18459 5069 18468
rect 4712 18284 4764 18290
rect 4540 18244 4712 18272
rect 4712 18226 4764 18232
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 4528 18148 4580 18154
rect 4528 18090 4580 18096
rect 4101 17980 4409 17989
rect 4101 17978 4107 17980
rect 4163 17978 4187 17980
rect 4243 17978 4267 17980
rect 4323 17978 4347 17980
rect 4403 17978 4409 17980
rect 4163 17926 4165 17978
rect 4345 17926 4347 17978
rect 4101 17924 4107 17926
rect 4163 17924 4187 17926
rect 4243 17924 4267 17926
rect 4323 17924 4347 17926
rect 4403 17924 4409 17926
rect 4101 17915 4409 17924
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4448 17202 4476 17682
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4101 16892 4409 16901
rect 4101 16890 4107 16892
rect 4163 16890 4187 16892
rect 4243 16890 4267 16892
rect 4323 16890 4347 16892
rect 4403 16890 4409 16892
rect 4163 16838 4165 16890
rect 4345 16838 4347 16890
rect 4101 16836 4107 16838
rect 4163 16836 4187 16838
rect 4243 16836 4267 16838
rect 4323 16836 4347 16838
rect 4403 16836 4409 16838
rect 4101 16827 4409 16836
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3804 15502 3832 16186
rect 3988 16046 4016 16390
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3896 15638 3924 15982
rect 4101 15804 4409 15813
rect 4101 15802 4107 15804
rect 4163 15802 4187 15804
rect 4243 15802 4267 15804
rect 4323 15802 4347 15804
rect 4403 15802 4409 15804
rect 4163 15750 4165 15802
rect 4345 15750 4347 15802
rect 4101 15748 4107 15750
rect 4163 15748 4187 15750
rect 4243 15748 4267 15750
rect 4323 15748 4347 15750
rect 4403 15748 4409 15750
rect 4101 15739 4409 15748
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 4540 15570 4568 18090
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4816 17882 4844 18022
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 5092 17746 5120 18158
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5184 17678 5212 18566
rect 5276 18426 5304 18634
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4712 17536 4764 17542
rect 4632 17496 4712 17524
rect 4632 16794 4660 17496
rect 4712 17478 4764 17484
rect 4761 17436 5069 17445
rect 4761 17434 4767 17436
rect 4823 17434 4847 17436
rect 4903 17434 4927 17436
rect 4983 17434 5007 17436
rect 5063 17434 5069 17436
rect 4823 17382 4825 17434
rect 5005 17382 5007 17434
rect 4761 17380 4767 17382
rect 4823 17380 4847 17382
rect 4903 17380 4927 17382
rect 4983 17380 5007 17382
rect 5063 17380 5069 17382
rect 4761 17371 5069 17380
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16794 4752 17070
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4761 16348 5069 16357
rect 4761 16346 4767 16348
rect 4823 16346 4847 16348
rect 4903 16346 4927 16348
rect 4983 16346 5007 16348
rect 5063 16346 5069 16348
rect 4823 16294 4825 16346
rect 5005 16294 5007 16346
rect 4761 16292 4767 16294
rect 4823 16292 4847 16294
rect 4903 16292 4927 16294
rect 4983 16292 5007 16294
rect 5063 16292 5069 16294
rect 4761 16283 5069 16292
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4540 14822 4568 15302
rect 4761 15260 5069 15269
rect 4761 15258 4767 15260
rect 4823 15258 4847 15260
rect 4903 15258 4927 15260
rect 4983 15258 5007 15260
rect 5063 15258 5069 15260
rect 4823 15206 4825 15258
rect 5005 15206 5007 15258
rect 4761 15204 4767 15206
rect 4823 15204 4847 15206
rect 4903 15204 4927 15206
rect 4983 15204 5007 15206
rect 5063 15204 5069 15206
rect 4761 15195 5069 15204
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4101 14716 4409 14725
rect 4101 14714 4107 14716
rect 4163 14714 4187 14716
rect 4243 14714 4267 14716
rect 4323 14714 4347 14716
rect 4403 14714 4409 14716
rect 4163 14662 4165 14714
rect 4345 14662 4347 14714
rect 4101 14660 4107 14662
rect 4163 14660 4187 14662
rect 4243 14660 4267 14662
rect 4323 14660 4347 14662
rect 4403 14660 4409 14662
rect 4101 14651 4409 14660
rect 4540 14414 4568 14758
rect 4908 14618 4936 14894
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 5184 14414 5212 15846
rect 5276 15502 5304 18362
rect 5368 18290 5396 19654
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5460 18222 5488 19858
rect 5644 19836 5672 21082
rect 5736 20398 5764 21966
rect 5920 21146 5948 21966
rect 5908 21140 5960 21146
rect 5960 21100 6040 21128
rect 5908 21082 5960 21088
rect 5816 20868 5868 20874
rect 5816 20810 5868 20816
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5736 20058 5764 20334
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5828 19854 5856 20810
rect 5920 20058 5948 20810
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 5724 19848 5776 19854
rect 5644 19808 5724 19836
rect 5724 19790 5776 19796
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5368 17678 5396 18022
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5368 16998 5396 17614
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5460 16182 5488 18022
rect 5552 17746 5580 18770
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5644 17542 5672 18090
rect 5736 17882 5764 19790
rect 5828 19378 5856 19790
rect 6012 19718 6040 21100
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6104 19854 6132 20198
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18290 6040 19110
rect 6196 18290 6224 22442
rect 6288 20466 6316 22578
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 21622 6684 21830
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6380 20534 6408 21422
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6368 20528 6420 20534
rect 6368 20470 6420 20476
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 6012 17678 6040 18226
rect 6288 17898 6316 20198
rect 6380 20074 6408 20470
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6380 20046 6500 20074
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6380 19378 6408 19926
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6380 18834 6408 19314
rect 6472 18970 6500 20046
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6104 17870 6316 17898
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5460 14958 5488 15982
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3804 12850 3832 13262
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3896 12238 3924 13806
rect 4101 13628 4409 13637
rect 4101 13626 4107 13628
rect 4163 13626 4187 13628
rect 4243 13626 4267 13628
rect 4323 13626 4347 13628
rect 4403 13626 4409 13628
rect 4163 13574 4165 13626
rect 4345 13574 4347 13626
rect 4101 13572 4107 13574
rect 4163 13572 4187 13574
rect 4243 13572 4267 13574
rect 4323 13572 4347 13574
rect 4403 13572 4409 13574
rect 4101 13563 4409 13572
rect 4448 12986 4476 13874
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4101 12540 4409 12549
rect 4101 12538 4107 12540
rect 4163 12538 4187 12540
rect 4243 12538 4267 12540
rect 4323 12538 4347 12540
rect 4403 12538 4409 12540
rect 4163 12486 4165 12538
rect 4345 12486 4347 12538
rect 4101 12484 4107 12486
rect 4163 12484 4187 12486
rect 4243 12484 4267 12486
rect 4323 12484 4347 12486
rect 4403 12484 4409 12486
rect 4101 12475 4409 12484
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 4342 12200 4398 12209
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11762 3832 12038
rect 3896 11812 3924 12174
rect 4342 12135 4344 12144
rect 4396 12135 4398 12144
rect 4344 12106 4396 12112
rect 4356 11898 4384 12106
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 3976 11824 4028 11830
rect 3896 11784 3976 11812
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3896 11626 3924 11784
rect 3976 11766 4028 11772
rect 4448 11626 4476 12786
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4101 11452 4409 11461
rect 4101 11450 4107 11452
rect 4163 11450 4187 11452
rect 4243 11450 4267 11452
rect 4323 11450 4347 11452
rect 4403 11450 4409 11452
rect 4163 11398 4165 11450
rect 4345 11398 4347 11450
rect 4101 11396 4107 11398
rect 4163 11396 4187 11398
rect 4243 11396 4267 11398
rect 4323 11396 4347 11398
rect 4403 11396 4409 11398
rect 4101 11387 4409 11396
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4101 10364 4409 10373
rect 4101 10362 4107 10364
rect 4163 10362 4187 10364
rect 4243 10362 4267 10364
rect 4323 10362 4347 10364
rect 4403 10362 4409 10364
rect 4163 10310 4165 10362
rect 4345 10310 4347 10362
rect 4101 10308 4107 10310
rect 4163 10308 4187 10310
rect 4243 10308 4267 10310
rect 4323 10308 4347 10310
rect 4403 10308 4409 10310
rect 4101 10299 4409 10308
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9586 3832 9862
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3804 8906 3832 9522
rect 4448 9382 4476 10950
rect 4540 10674 4568 14350
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4632 14006 4660 14214
rect 4761 14172 5069 14181
rect 4761 14170 4767 14172
rect 4823 14170 4847 14172
rect 4903 14170 4927 14172
rect 4983 14170 5007 14172
rect 5063 14170 5069 14172
rect 4823 14118 4825 14170
rect 5005 14118 5007 14170
rect 4761 14116 4767 14118
rect 4823 14116 4847 14118
rect 4903 14116 4927 14118
rect 4983 14116 5007 14118
rect 5063 14116 5069 14118
rect 4761 14107 5069 14116
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 11354 4660 13670
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 4761 13084 5069 13093
rect 4761 13082 4767 13084
rect 4823 13082 4847 13084
rect 4903 13082 4927 13084
rect 4983 13082 5007 13084
rect 5063 13082 5069 13084
rect 4823 13030 4825 13082
rect 5005 13030 5007 13082
rect 4761 13028 4767 13030
rect 4823 13028 4847 13030
rect 4903 13028 4927 13030
rect 4983 13028 5007 13030
rect 5063 13028 5069 13030
rect 4761 13019 5069 13028
rect 5184 12986 5212 13262
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4816 12374 4844 12922
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 5184 12238 5212 12922
rect 5276 12850 5304 13398
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 4761 11996 5069 12005
rect 4761 11994 4767 11996
rect 4823 11994 4847 11996
rect 4903 11994 4927 11996
rect 4983 11994 5007 11996
rect 5063 11994 5069 11996
rect 4823 11942 4825 11994
rect 5005 11942 5007 11994
rect 4761 11940 4767 11942
rect 4823 11940 4847 11942
rect 4903 11940 4927 11942
rect 4983 11940 5007 11942
rect 5063 11940 5069 11942
rect 4761 11931 5069 11940
rect 4710 11792 4766 11801
rect 4710 11727 4712 11736
rect 4764 11727 4766 11736
rect 4896 11756 4948 11762
rect 4712 11698 4764 11704
rect 4896 11698 4948 11704
rect 4908 11354 4936 11698
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5184 11218 5212 12174
rect 5276 11286 5304 12650
rect 5460 12345 5488 14894
rect 5552 14346 5580 16390
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5446 12336 5502 12345
rect 5552 12306 5580 12582
rect 5644 12434 5672 17478
rect 6012 17202 6040 17478
rect 6000 17196 6052 17202
rect 5828 17156 6000 17184
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5736 16590 5764 17002
rect 5828 16658 5856 17156
rect 6000 17138 6052 17144
rect 6104 16946 6132 17870
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6196 17542 6224 17750
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6012 16918 6132 16946
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 6012 15910 6040 16918
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6104 16590 6132 16730
rect 6196 16590 6224 17206
rect 6288 16658 6316 17478
rect 6380 16998 6408 18770
rect 6564 18766 6592 20402
rect 6656 19990 6684 20946
rect 6748 20806 6776 21966
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 21622 7144 21830
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6748 20398 6776 20742
rect 6932 20602 6960 21082
rect 7484 21078 7512 21898
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 7472 21072 7524 21078
rect 7472 21014 7524 21020
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6748 20262 6776 20334
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6472 17270 6500 17818
rect 6656 17678 6684 19722
rect 6736 19712 6788 19718
rect 6840 19700 6868 20334
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6788 19672 6868 19700
rect 6736 19654 6788 19660
rect 6748 19378 6776 19654
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6748 17882 6776 19314
rect 6828 18216 6880 18222
rect 6932 18170 6960 19994
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7116 18766 7144 19858
rect 7300 19854 7328 21014
rect 7484 20602 7512 21014
rect 7668 20942 7696 21286
rect 8036 21146 8064 21354
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8680 20942 8708 21490
rect 8772 21146 8800 21966
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8956 21622 8984 21830
rect 9140 21690 9168 21966
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 7656 20936 7708 20942
rect 8668 20936 8720 20942
rect 7656 20878 7708 20884
rect 8588 20896 8668 20924
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7668 19922 7696 20878
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7208 18970 7236 19382
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 6880 18164 6960 18170
rect 6828 18158 6960 18164
rect 6840 18142 6960 18158
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6644 17536 6696 17542
rect 6642 17504 6644 17513
rect 6696 17504 6698 17513
rect 6642 17439 6698 17448
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6472 16726 6500 17206
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6460 16720 6512 16726
rect 6460 16662 6512 16668
rect 6564 16658 6592 17070
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6012 15706 6040 15846
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5736 14618 5764 15030
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 6012 14414 6040 15642
rect 6380 14414 6408 15846
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6472 14362 6500 15574
rect 6564 15366 6592 16594
rect 6656 16454 6684 17439
rect 6748 17082 6776 17818
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17202 6868 17614
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6932 17116 6960 18142
rect 7104 17672 7156 17678
rect 7208 17660 7236 18906
rect 7944 17921 7972 19722
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 8036 19378 8064 19654
rect 8496 19514 8524 20334
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8588 18426 8616 20896
rect 8668 20878 8720 20884
rect 9232 20618 9260 22646
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9324 21486 9352 21966
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 9140 20590 9260 20618
rect 9324 20602 9352 21422
rect 9416 21010 9444 22646
rect 10796 22630 10916 22658
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 9784 21350 9812 22374
rect 10336 21962 10364 22374
rect 10403 22332 10711 22341
rect 10403 22330 10409 22332
rect 10465 22330 10489 22332
rect 10545 22330 10569 22332
rect 10625 22330 10649 22332
rect 10705 22330 10711 22332
rect 10465 22278 10467 22330
rect 10647 22278 10649 22330
rect 10403 22276 10409 22278
rect 10465 22276 10489 22278
rect 10545 22276 10569 22278
rect 10625 22276 10649 22278
rect 10705 22276 10711 22278
rect 10403 22267 10711 22276
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 10403 21244 10711 21253
rect 10403 21242 10409 21244
rect 10465 21242 10489 21244
rect 10545 21242 10569 21244
rect 10625 21242 10649 21244
rect 10705 21242 10711 21244
rect 10465 21190 10467 21242
rect 10647 21190 10649 21242
rect 10403 21188 10409 21190
rect 10465 21188 10489 21190
rect 10545 21188 10569 21190
rect 10625 21188 10649 21190
rect 10705 21188 10711 21190
rect 10403 21179 10711 21188
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 10796 20602 10824 22630
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 10888 21622 10916 22374
rect 11348 22234 11376 22374
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11063 21788 11371 21797
rect 11063 21786 11069 21788
rect 11125 21786 11149 21788
rect 11205 21786 11229 21788
rect 11285 21786 11309 21788
rect 11365 21786 11371 21788
rect 11125 21734 11127 21786
rect 11307 21734 11309 21786
rect 11063 21732 11069 21734
rect 11125 21732 11149 21734
rect 11205 21732 11229 21734
rect 11285 21732 11309 21734
rect 11365 21732 11371 21734
rect 11063 21723 11371 21732
rect 10876 21616 10928 21622
rect 10876 21558 10928 21564
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 9312 20596 9364 20602
rect 9140 19854 9168 20590
rect 9312 20538 9364 20544
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 9232 20058 9260 20470
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9324 19922 9352 20538
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 7930 17912 7986 17921
rect 7472 17876 7524 17882
rect 7930 17847 7986 17856
rect 7472 17818 7524 17824
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7156 17632 7236 17660
rect 7104 17614 7156 17620
rect 7208 17592 7236 17632
rect 7288 17604 7340 17610
rect 7208 17564 7288 17592
rect 7288 17546 7340 17552
rect 7012 17128 7064 17134
rect 6932 17088 7012 17116
rect 6748 17054 6868 17082
rect 7012 17070 7064 17076
rect 6840 16998 6868 17054
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6656 16250 6684 16390
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6748 15978 6776 16934
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 15162 6592 15302
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6564 14550 6592 15098
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6656 14618 6684 14894
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6472 14334 6592 14362
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5920 13938 5948 14214
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 5920 13530 5948 13670
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5644 12406 5764 12434
rect 5630 12336 5686 12345
rect 5446 12271 5502 12280
rect 5540 12300 5592 12306
rect 5630 12271 5686 12280
rect 5540 12242 5592 12248
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11801 5396 12038
rect 5354 11792 5410 11801
rect 5354 11727 5410 11736
rect 5460 11354 5488 12174
rect 5540 11824 5592 11830
rect 5538 11792 5540 11801
rect 5592 11792 5594 11801
rect 5644 11762 5672 12271
rect 5538 11727 5594 11736
rect 5637 11756 5689 11762
rect 5637 11698 5689 11704
rect 5644 11665 5672 11698
rect 5630 11656 5686 11665
rect 5630 11591 5686 11600
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5736 11286 5764 12406
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5828 11898 5856 12106
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5920 11558 5948 13466
rect 6104 13394 6132 13670
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6196 12442 6224 13262
rect 6564 12782 6592 14334
rect 6748 14278 6776 14894
rect 6840 14414 6868 16730
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7300 16250 7328 16458
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7392 15570 7420 17750
rect 7484 17338 7512 17818
rect 7944 17542 7972 17847
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 8404 16114 8432 17750
rect 8588 16182 8616 18362
rect 8772 18222 8800 18566
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8680 16794 8708 17478
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 7116 14618 7144 15030
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13954 6776 14214
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6656 13926 6776 13954
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6184 12436 6236 12442
rect 6564 12434 6592 12718
rect 6184 12378 6236 12384
rect 6472 12406 6592 12434
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11778 6040 12038
rect 6104 11898 6132 12174
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6012 11762 6132 11778
rect 6012 11756 6144 11762
rect 6012 11750 6092 11756
rect 6092 11698 6144 11704
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 6012 11354 6040 11630
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5264 11280 5316 11286
rect 5540 11280 5592 11286
rect 5264 11222 5316 11228
rect 5538 11248 5540 11257
rect 5724 11280 5776 11286
rect 5592 11248 5594 11257
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5276 11014 5304 11222
rect 5724 11222 5776 11228
rect 5538 11183 5594 11192
rect 6104 11014 6132 11698
rect 6196 11150 6224 12378
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11830 6316 12174
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6288 11354 6316 11562
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6368 11280 6420 11286
rect 6366 11248 6368 11257
rect 6420 11248 6422 11257
rect 6276 11212 6328 11218
rect 6366 11183 6422 11192
rect 6276 11154 6328 11160
rect 6184 11144 6236 11150
rect 6288 11121 6316 11154
rect 6184 11086 6236 11092
rect 6274 11112 6330 11121
rect 6472 11082 6500 12406
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6564 11150 6592 12242
rect 6656 12238 6684 13926
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13530 6776 13738
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6748 12714 6776 13466
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6644 12232 6696 12238
rect 6840 12209 6868 14010
rect 7300 13938 7328 15302
rect 7576 15162 7604 15982
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7944 15502 7972 15642
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8128 15162 8156 15438
rect 8588 15434 8616 16118
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7392 14074 7420 14282
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7668 14006 7696 14826
rect 8312 14346 8340 15302
rect 8588 15094 8616 15370
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 14006 8708 14214
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7024 13530 7052 13874
rect 7208 13818 7236 13874
rect 7208 13790 7328 13818
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6644 12174 6696 12180
rect 6826 12200 6882 12209
rect 6656 11898 6684 12174
rect 6882 12158 6960 12186
rect 6826 12135 6882 12144
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6734 11792 6790 11801
rect 6734 11727 6736 11736
rect 6788 11727 6790 11736
rect 6736 11698 6788 11704
rect 6734 11656 6790 11665
rect 6734 11591 6790 11600
rect 6748 11558 6776 11591
rect 6736 11552 6788 11558
rect 6656 11512 6736 11540
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6274 11047 6330 11056
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 4761 10908 5069 10917
rect 4761 10906 4767 10908
rect 4823 10906 4847 10908
rect 4903 10906 4927 10908
rect 4983 10906 5007 10908
rect 5063 10906 5069 10908
rect 4823 10854 4825 10906
rect 5005 10854 5007 10906
rect 4761 10852 4767 10854
rect 4823 10852 4847 10854
rect 4903 10852 4927 10854
rect 4983 10852 5007 10854
rect 5063 10852 5069 10854
rect 4761 10843 5069 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4632 9674 4660 10610
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5184 10062 5212 10474
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 4761 9820 5069 9829
rect 4761 9818 4767 9820
rect 4823 9818 4847 9820
rect 4903 9818 4927 9820
rect 4983 9818 5007 9820
rect 5063 9818 5069 9820
rect 4823 9766 4825 9818
rect 5005 9766 5007 9818
rect 4761 9764 4767 9766
rect 4823 9764 4847 9766
rect 4903 9764 4927 9766
rect 4983 9764 5007 9766
rect 5063 9764 5069 9766
rect 4761 9755 5069 9764
rect 4632 9646 5028 9674
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4101 9276 4409 9285
rect 4101 9274 4107 9276
rect 4163 9274 4187 9276
rect 4243 9274 4267 9276
rect 4323 9274 4347 9276
rect 4403 9274 4409 9276
rect 4163 9222 4165 9274
rect 4345 9222 4347 9274
rect 4101 9220 4107 9222
rect 4163 9220 4187 9222
rect 4243 9220 4267 9222
rect 4323 9220 4347 9222
rect 4403 9220 4409 9222
rect 4101 9211 4409 9220
rect 4448 9110 4476 9318
rect 4632 9178 4660 9522
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4436 9104 4488 9110
rect 4804 9104 4856 9110
rect 4436 9046 4488 9052
rect 4802 9072 4804 9081
rect 4856 9072 4858 9081
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 4172 8634 4200 9046
rect 4802 9007 4858 9016
rect 4620 8968 4672 8974
rect 4908 8945 4936 9522
rect 5000 8956 5028 9646
rect 5184 9568 5212 9998
rect 5092 9540 5212 9568
rect 5092 9382 5120 9540
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5172 8968 5224 8974
rect 4620 8910 4672 8916
rect 4894 8936 4950 8945
rect 4632 8650 4660 8910
rect 5000 8928 5172 8956
rect 5172 8910 5224 8916
rect 4894 8871 4950 8880
rect 4761 8732 5069 8741
rect 4761 8730 4767 8732
rect 4823 8730 4847 8732
rect 4903 8730 4927 8732
rect 4983 8730 5007 8732
rect 5063 8730 5069 8732
rect 4823 8678 4825 8730
rect 5005 8678 5007 8730
rect 4761 8676 4767 8678
rect 4823 8676 4847 8678
rect 4903 8676 4927 8678
rect 4983 8676 5007 8678
rect 5063 8676 5069 8678
rect 4761 8667 5069 8676
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4448 8622 4660 8650
rect 4101 8188 4409 8197
rect 4101 8186 4107 8188
rect 4163 8186 4187 8188
rect 4243 8186 4267 8188
rect 4323 8186 4347 8188
rect 4403 8186 4409 8188
rect 4163 8134 4165 8186
rect 4345 8134 4347 8186
rect 4101 8132 4107 8134
rect 4163 8132 4187 8134
rect 4243 8132 4267 8134
rect 4323 8132 4347 8134
rect 4403 8132 4409 8134
rect 4101 8123 4409 8132
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4172 7410 4200 7822
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4264 7324 4292 7822
rect 4448 7818 4476 8622
rect 4632 8566 4660 8622
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4620 8560 4672 8566
rect 5000 8537 5028 8570
rect 4620 8502 4672 8508
rect 4986 8528 5042 8537
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4448 7546 4476 7754
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4344 7336 4396 7342
rect 4264 7296 4344 7324
rect 4344 7278 4396 7284
rect 4540 7274 4568 8502
rect 4986 8463 5042 8472
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 7410 4660 8230
rect 4724 8022 4752 8298
rect 4712 8016 4764 8022
rect 5184 7970 5212 8910
rect 4712 7958 4764 7964
rect 5092 7942 5212 7970
rect 5092 7818 5120 7942
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4761 7644 5069 7653
rect 4761 7642 4767 7644
rect 4823 7642 4847 7644
rect 4903 7642 4927 7644
rect 4983 7642 5007 7644
rect 5063 7642 5069 7644
rect 4823 7590 4825 7642
rect 5005 7590 5007 7642
rect 4761 7588 4767 7590
rect 4823 7588 4847 7590
rect 4903 7588 4927 7590
rect 4983 7588 5007 7590
rect 5063 7588 5069 7590
rect 4761 7579 5069 7588
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 3804 6798 3832 7142
rect 4101 7100 4409 7109
rect 4101 7098 4107 7100
rect 4163 7098 4187 7100
rect 4243 7098 4267 7100
rect 4323 7098 4347 7100
rect 4403 7098 4409 7100
rect 4163 7046 4165 7098
rect 4345 7046 4347 7098
rect 4101 7044 4107 7046
rect 4163 7044 4187 7046
rect 4243 7044 4267 7046
rect 4323 7044 4347 7046
rect 4403 7044 4409 7046
rect 4101 7035 4409 7044
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 5914 3832 6734
rect 4724 6730 4752 7142
rect 5184 7002 5212 7822
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4761 6556 5069 6565
rect 4761 6554 4767 6556
rect 4823 6554 4847 6556
rect 4903 6554 4927 6556
rect 4983 6554 5007 6556
rect 5063 6554 5069 6556
rect 4823 6502 4825 6554
rect 5005 6502 5007 6554
rect 4761 6500 4767 6502
rect 4823 6500 4847 6502
rect 4903 6500 4927 6502
rect 4983 6500 5007 6502
rect 5063 6500 5069 6502
rect 4761 6491 5069 6500
rect 4101 6012 4409 6021
rect 4101 6010 4107 6012
rect 4163 6010 4187 6012
rect 4243 6010 4267 6012
rect 4323 6010 4347 6012
rect 4403 6010 4409 6012
rect 4163 5958 4165 6010
rect 4345 5958 4347 6010
rect 4101 5956 4107 5958
rect 4163 5956 4187 5958
rect 4243 5956 4267 5958
rect 4323 5956 4347 5958
rect 4403 5956 4409 5958
rect 4101 5947 4409 5956
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 5276 5710 5304 9998
rect 5368 6186 5396 10406
rect 5460 9518 5488 10746
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5552 8838 5580 10542
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 9654 5672 10406
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5538 8664 5594 8673
rect 5448 8628 5500 8634
rect 5538 8599 5594 8608
rect 5448 8570 5500 8576
rect 5460 7002 5488 8570
rect 5552 8498 5580 8599
rect 5644 8498 5672 9046
rect 5828 8974 5856 9318
rect 5920 9042 5948 9998
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6012 9654 6040 9930
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6104 9586 6132 10950
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5724 8964 5776 8970
rect 5724 8906 5776 8912
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 6012 8906 6040 8978
rect 5736 8634 5764 8906
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5724 8628 5776 8634
rect 6012 8616 6040 8842
rect 5724 8570 5776 8576
rect 5828 8588 6040 8616
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5552 7868 5580 8434
rect 5828 8362 5856 8588
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5630 8120 5686 8129
rect 5630 8055 5686 8064
rect 5644 8022 5672 8055
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5920 7954 5948 8434
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5552 7840 5672 7868
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5552 6458 5580 6734
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4761 5468 5069 5477
rect 4761 5466 4767 5468
rect 4823 5466 4847 5468
rect 4903 5466 4927 5468
rect 4983 5466 5007 5468
rect 5063 5466 5069 5468
rect 4823 5414 4825 5466
rect 5005 5414 5007 5466
rect 4761 5412 4767 5414
rect 4823 5412 4847 5414
rect 4903 5412 4927 5414
rect 4983 5412 5007 5414
rect 5063 5412 5069 5414
rect 4761 5403 5069 5412
rect 4101 4924 4409 4933
rect 4101 4922 4107 4924
rect 4163 4922 4187 4924
rect 4243 4922 4267 4924
rect 4323 4922 4347 4924
rect 4403 4922 4409 4924
rect 4163 4870 4165 4922
rect 4345 4870 4347 4922
rect 4101 4868 4107 4870
rect 4163 4868 4187 4870
rect 4243 4868 4267 4870
rect 4323 4868 4347 4870
rect 4403 4868 4409 4870
rect 4101 4859 4409 4868
rect 5552 4622 5580 6394
rect 5644 6186 5672 7840
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5736 5370 5764 6258
rect 6012 5710 6040 8588
rect 6104 6322 6132 9522
rect 6288 9382 6316 10678
rect 6564 9926 6592 11086
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 8838 6316 9318
rect 6380 8974 6408 9862
rect 6564 9722 6592 9862
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6458 9072 6514 9081
rect 6458 9007 6460 9016
rect 6512 9007 6514 9016
rect 6460 8978 6512 8984
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6552 8900 6604 8906
rect 6656 8888 6684 11512
rect 6736 11494 6788 11500
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6748 8906 6776 10202
rect 6840 9994 6868 12038
rect 6932 10266 6960 12158
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6840 9178 6868 9930
rect 7024 9674 7052 12582
rect 7208 11694 7236 13330
rect 7300 13190 7328 13790
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12442 7328 13126
rect 7392 12850 7420 13670
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7484 12730 7512 13942
rect 8772 13802 8800 17478
rect 8956 17202 8984 17478
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9048 17134 9076 18022
rect 9140 17678 9168 19790
rect 9324 19446 9352 19858
rect 9600 19854 9628 20266
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9968 20058 9996 20198
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9508 19258 9536 19314
rect 9508 19230 9720 19258
rect 9692 18970 9720 19230
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8956 14958 8984 16934
rect 9140 16726 9168 17614
rect 9324 17338 9352 18294
rect 9968 18222 9996 19994
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9324 17134 9352 17274
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9140 16590 9168 16662
rect 9784 16590 9812 17206
rect 9968 17066 9996 18158
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 10060 16726 10088 20538
rect 10980 20534 11008 20810
rect 11063 20700 11371 20709
rect 11063 20698 11069 20700
rect 11125 20698 11149 20700
rect 11205 20698 11229 20700
rect 11285 20698 11309 20700
rect 11365 20698 11371 20700
rect 11125 20646 11127 20698
rect 11307 20646 11309 20698
rect 11063 20644 11069 20646
rect 11125 20644 11149 20646
rect 11205 20644 11229 20646
rect 11285 20644 11309 20646
rect 11365 20644 11371 20646
rect 11063 20635 11371 20644
rect 10140 20528 10192 20534
rect 10140 20470 10192 20476
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10152 18630 10180 20470
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 10403 20156 10711 20165
rect 10403 20154 10409 20156
rect 10465 20154 10489 20156
rect 10545 20154 10569 20156
rect 10625 20154 10649 20156
rect 10705 20154 10711 20156
rect 10465 20102 10467 20154
rect 10647 20102 10649 20154
rect 10403 20100 10409 20102
rect 10465 20100 10489 20102
rect 10545 20100 10569 20102
rect 10625 20100 10649 20102
rect 10705 20100 10711 20102
rect 10403 20091 10711 20100
rect 11440 20058 11468 20402
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11063 19612 11371 19621
rect 11063 19610 11069 19612
rect 11125 19610 11149 19612
rect 11205 19610 11229 19612
rect 11285 19610 11309 19612
rect 11365 19610 11371 19612
rect 11125 19558 11127 19610
rect 11307 19558 11309 19610
rect 11063 19556 11069 19558
rect 11125 19556 11149 19558
rect 11205 19556 11229 19558
rect 11285 19556 11309 19558
rect 11365 19556 11371 19558
rect 11063 19547 11371 19556
rect 10322 19408 10378 19417
rect 10322 19343 10378 19352
rect 10336 18834 10364 19343
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 10403 19068 10711 19077
rect 10403 19066 10409 19068
rect 10465 19066 10489 19068
rect 10545 19066 10569 19068
rect 10625 19066 10649 19068
rect 10705 19066 10711 19068
rect 10465 19014 10467 19066
rect 10647 19014 10649 19066
rect 10403 19012 10409 19014
rect 10465 19012 10489 19014
rect 10545 19012 10569 19014
rect 10625 19012 10649 19014
rect 10705 19012 10711 19014
rect 10403 19003 10711 19012
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 11348 18698 11376 19110
rect 11440 18970 11468 19790
rect 11532 19496 11560 26930
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11900 25906 11928 26318
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11612 25696 11664 25702
rect 11612 25638 11664 25644
rect 11624 25294 11652 25638
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11900 24206 11928 25842
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11624 23866 11652 24142
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11716 22778 11744 23462
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 11624 21894 11652 22578
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11624 21010 11652 21830
rect 11900 21146 11928 24142
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 23662 12112 24006
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11992 22778 12020 22918
rect 12084 22778 12112 23598
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11992 22166 12020 22578
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11992 22030 12020 22102
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12084 21554 12112 21966
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11532 19468 11652 19496
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11532 18766 11560 19314
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10152 17921 10180 18566
rect 11063 18524 11371 18533
rect 11063 18522 11069 18524
rect 11125 18522 11149 18524
rect 11205 18522 11229 18524
rect 11285 18522 11309 18524
rect 11365 18522 11371 18524
rect 11125 18470 11127 18522
rect 11307 18470 11309 18522
rect 11063 18468 11069 18470
rect 11125 18468 11149 18470
rect 11205 18468 11229 18470
rect 11285 18468 11309 18470
rect 11365 18468 11371 18470
rect 11063 18459 11371 18468
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10138 17912 10194 17921
rect 10138 17847 10194 17856
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10152 17338 10180 17546
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10244 16998 10272 17750
rect 10336 17202 10364 18294
rect 10796 18290 10824 18362
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10403 17980 10711 17989
rect 10403 17978 10409 17980
rect 10465 17978 10489 17980
rect 10545 17978 10569 17980
rect 10625 17978 10649 17980
rect 10705 17978 10711 17980
rect 10465 17926 10467 17978
rect 10647 17926 10649 17978
rect 10403 17924 10409 17926
rect 10465 17924 10489 17926
rect 10545 17924 10569 17926
rect 10625 17924 10649 17926
rect 10705 17924 10711 17926
rect 10403 17915 10711 17924
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9784 16114 9812 16526
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9968 15502 9996 16662
rect 10244 16504 10272 16934
rect 10336 16658 10364 17138
rect 10403 16892 10711 16901
rect 10403 16890 10409 16892
rect 10465 16890 10489 16892
rect 10545 16890 10569 16892
rect 10625 16890 10649 16892
rect 10705 16890 10711 16892
rect 10465 16838 10467 16890
rect 10647 16838 10649 16890
rect 10403 16836 10409 16838
rect 10465 16836 10489 16838
rect 10545 16836 10569 16838
rect 10625 16836 10649 16838
rect 10705 16836 10711 16838
rect 10403 16827 10711 16836
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10324 16516 10376 16522
rect 10244 16476 10324 16504
rect 10324 16458 10376 16464
rect 10336 16250 10364 16458
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10796 16114 10824 18022
rect 10888 17814 10916 18226
rect 11072 18170 11100 18226
rect 11072 18142 11376 18170
rect 11348 18086 11376 18142
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 11520 17604 11572 17610
rect 11520 17546 11572 17552
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11063 17436 11371 17445
rect 11063 17434 11069 17436
rect 11125 17434 11149 17436
rect 11205 17434 11229 17436
rect 11285 17434 11309 17436
rect 11365 17434 11371 17436
rect 11125 17382 11127 17434
rect 11307 17382 11309 17434
rect 11063 17380 11069 17382
rect 11125 17380 11149 17382
rect 11205 17380 11229 17382
rect 11285 17380 11309 17382
rect 11365 17380 11371 17382
rect 11063 17371 11371 17380
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10888 16998 10916 17138
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10888 16046 10916 16934
rect 11440 16658 11468 17478
rect 11532 17338 11560 17546
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11624 17202 11652 19468
rect 11716 18290 11744 19994
rect 12084 19446 12112 21490
rect 12360 20058 12388 26930
rect 16304 26784 16356 26790
rect 16304 26726 16356 26732
rect 13728 26444 13780 26450
rect 13728 26386 13780 26392
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12452 25430 12480 26318
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 12716 25968 12768 25974
rect 12716 25910 12768 25916
rect 12728 25498 12756 25910
rect 12820 25498 12848 25978
rect 13740 25906 13768 26386
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 13832 26042 13860 26318
rect 15476 26308 15528 26314
rect 15476 26250 15528 26256
rect 14648 26240 14700 26246
rect 14648 26182 14700 26188
rect 14660 26042 14688 26182
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 13728 25900 13780 25906
rect 13728 25842 13780 25848
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 12716 25492 12768 25498
rect 12716 25434 12768 25440
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12440 25424 12492 25430
rect 12440 25366 12492 25372
rect 12820 25294 12848 25434
rect 13084 25424 13136 25430
rect 13084 25366 13136 25372
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 13096 24954 13124 25366
rect 13084 24948 13136 24954
rect 13084 24890 13136 24896
rect 13464 24682 13492 25638
rect 13740 25498 13768 25842
rect 14004 25696 14056 25702
rect 14004 25638 14056 25644
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13544 25424 13596 25430
rect 13544 25366 13596 25372
rect 13556 24886 13584 25366
rect 13544 24880 13596 24886
rect 13544 24822 13596 24828
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13452 24676 13504 24682
rect 13452 24618 13504 24624
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12452 24274 12480 24550
rect 13648 24274 13676 24754
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 13636 24268 13688 24274
rect 13636 24210 13688 24216
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23866 13032 24074
rect 13648 23866 13676 24210
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13740 23730 13768 25434
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13832 24954 13860 25230
rect 13820 24948 13872 24954
rect 13820 24890 13872 24896
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 13832 23730 13860 24142
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 12820 22574 12848 23530
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 21690 12480 22374
rect 12544 21894 12572 22510
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12716 22094 12768 22098
rect 12820 22094 12848 22374
rect 12716 22092 12848 22094
rect 12768 22066 12848 22092
rect 12716 22034 12768 22040
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12912 20942 12940 23666
rect 13924 23662 13952 24754
rect 14016 24206 14044 25638
rect 14660 25294 14688 25978
rect 15488 25974 15516 26250
rect 15948 26042 15976 26318
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 15476 25968 15528 25974
rect 15476 25910 15528 25916
rect 16316 25906 16344 26726
rect 16705 26684 17013 26693
rect 16705 26682 16711 26684
rect 16767 26682 16791 26684
rect 16847 26682 16871 26684
rect 16927 26682 16951 26684
rect 17007 26682 17013 26684
rect 16767 26630 16769 26682
rect 16949 26630 16951 26682
rect 16705 26628 16711 26630
rect 16767 26628 16791 26630
rect 16847 26628 16871 26630
rect 16927 26628 16951 26630
rect 17007 26628 17013 26630
rect 16705 26619 17013 26628
rect 18420 26444 18472 26450
rect 18420 26386 18472 26392
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 16304 25900 16356 25906
rect 16304 25842 16356 25848
rect 15476 25832 15528 25838
rect 15476 25774 15528 25780
rect 15488 25498 15516 25774
rect 15844 25764 15896 25770
rect 15844 25706 15896 25712
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24886 14412 25094
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 14844 24818 14872 25298
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15752 25288 15804 25294
rect 15752 25230 15804 25236
rect 14936 25158 14964 25230
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14936 24954 14964 25094
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 13004 22778 13032 23122
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 13004 22098 13032 22510
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 13740 22012 13768 22374
rect 14292 22030 14320 23666
rect 14476 23594 14504 24754
rect 14660 24410 14688 24754
rect 14936 24682 14964 24890
rect 15028 24886 15056 25162
rect 15304 24954 15332 25230
rect 15764 24954 15792 25230
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 15212 24410 15240 24754
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15764 24410 15792 24686
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 14660 23730 14688 24210
rect 14752 24206 14780 24278
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14936 23798 14964 24346
rect 15660 24268 15712 24274
rect 15660 24210 15712 24216
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 15304 23798 15332 24074
rect 15580 23798 15608 24142
rect 15672 24120 15700 24210
rect 15752 24132 15804 24138
rect 15672 24092 15752 24120
rect 14924 23792 14976 23798
rect 14924 23734 14976 23740
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 15672 23662 15700 24092
rect 15752 24074 15804 24080
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 14464 23588 14516 23594
rect 14464 23530 14516 23536
rect 15672 22710 15700 23598
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15028 22098 15056 22578
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 13912 22024 13964 22030
rect 13740 21984 13912 22012
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 13096 21146 13124 21898
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13648 21350 13676 21830
rect 13740 21690 13768 21984
rect 13912 21966 13964 21972
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 14108 21078 14136 21422
rect 14292 21418 14320 21966
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14372 21616 14424 21622
rect 14372 21558 14424 21564
rect 14280 21412 14332 21418
rect 14280 21354 14332 21360
rect 14384 21146 14412 21558
rect 14476 21554 14504 21830
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 13268 20936 13320 20942
rect 14280 20936 14332 20942
rect 13268 20878 13320 20884
rect 14278 20904 14280 20913
rect 14332 20904 14334 20913
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11900 18290 11928 18362
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11348 16504 11376 16594
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11348 16476 11468 16504
rect 11063 16348 11371 16357
rect 11063 16346 11069 16348
rect 11125 16346 11149 16348
rect 11205 16346 11229 16348
rect 11285 16346 11309 16348
rect 11365 16346 11371 16348
rect 11125 16294 11127 16346
rect 11307 16294 11309 16346
rect 11063 16292 11069 16294
rect 11125 16292 11149 16294
rect 11205 16292 11229 16294
rect 11285 16292 11309 16294
rect 11365 16292 11371 16294
rect 11063 16283 11371 16292
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10403 15804 10711 15813
rect 10403 15802 10409 15804
rect 10465 15802 10489 15804
rect 10545 15802 10569 15804
rect 10625 15802 10649 15804
rect 10705 15802 10711 15804
rect 10465 15750 10467 15802
rect 10647 15750 10649 15802
rect 10403 15748 10409 15750
rect 10465 15748 10489 15750
rect 10545 15748 10569 15750
rect 10625 15748 10649 15750
rect 10705 15748 10711 15750
rect 10403 15739 10711 15748
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7392 12702 7512 12730
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7392 11830 7420 12702
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7484 11762 7512 12582
rect 7668 12102 7696 13262
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7668 11694 7696 12038
rect 8128 11830 8156 12718
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 12209 8248 12242
rect 8312 12238 8340 12582
rect 8300 12232 8352 12238
rect 8206 12200 8262 12209
rect 8300 12174 8352 12180
rect 8206 12135 8262 12144
rect 8404 11898 8432 12650
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7208 11218 7236 11630
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7668 11121 7696 11630
rect 7654 11112 7710 11121
rect 8496 11082 8524 12310
rect 8588 12238 8616 12786
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 11354 8616 11630
rect 8864 11354 8892 14894
rect 9232 14482 9260 14894
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9140 14074 9168 14350
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9324 13938 9352 15302
rect 9784 15094 9812 15302
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9876 14822 9904 15438
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10152 15094 10180 15302
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 10244 14346 10272 15302
rect 11063 15260 11371 15269
rect 11063 15258 11069 15260
rect 11125 15258 11149 15260
rect 11205 15258 11229 15260
rect 11285 15258 11309 15260
rect 11365 15258 11371 15260
rect 11125 15206 11127 15258
rect 11307 15206 11309 15258
rect 11063 15204 11069 15206
rect 11125 15204 11149 15206
rect 11205 15204 11229 15206
rect 11285 15204 11309 15206
rect 11365 15204 11371 15206
rect 11063 15195 11371 15204
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10403 14716 10711 14725
rect 10403 14714 10409 14716
rect 10465 14714 10489 14716
rect 10545 14714 10569 14716
rect 10625 14714 10649 14716
rect 10705 14714 10711 14716
rect 10465 14662 10467 14714
rect 10647 14662 10649 14714
rect 10403 14660 10409 14662
rect 10465 14660 10489 14662
rect 10545 14660 10569 14662
rect 10625 14660 10649 14662
rect 10705 14660 10711 14662
rect 10403 14651 10711 14660
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9508 13870 9536 14010
rect 10796 14006 10824 14962
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9508 12850 9536 13806
rect 9692 12974 9996 13002
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 7654 11047 7710 11056
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8588 10606 8616 11290
rect 8956 10674 8984 12718
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9232 11694 9260 12106
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9232 11150 9260 11630
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9324 10810 9352 12174
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9508 10674 9536 12786
rect 9692 12714 9720 12974
rect 9968 12918 9996 12974
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 10060 12850 10088 13942
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11762 9628 12038
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9784 11218 9812 12650
rect 9876 11642 9904 12786
rect 10060 11694 10088 12786
rect 10152 11898 10180 12786
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11688 10100 11694
rect 9876 11614 9996 11642
rect 10048 11630 10100 11636
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9968 11082 9996 11614
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8956 10266 8984 10610
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9692 10062 9720 10542
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 6932 9646 7052 9674
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6604 8860 6684 8888
rect 6736 8900 6788 8906
rect 6552 8842 6604 8848
rect 6736 8842 6788 8848
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6288 8090 6316 8502
rect 6840 8362 6868 9114
rect 6932 8634 6960 9646
rect 7576 9586 7604 9862
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9178 8064 9522
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6932 8242 6960 8570
rect 8128 8498 8156 8978
rect 9140 8974 9168 9998
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 6748 8214 6960 8242
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6380 7002 6408 7958
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 6322 6592 6598
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6104 5642 6132 6258
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 6196 5846 6224 6122
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 6656 5234 6684 6394
rect 6748 5302 6776 8214
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 7002 7512 7142
rect 7668 7002 7696 7822
rect 8128 7410 8156 8434
rect 8404 8090 8432 8434
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6840 6322 6868 6394
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6656 4842 6684 5170
rect 6840 5166 6868 5646
rect 6932 5234 6960 6598
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 7024 5030 7052 6802
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7116 5778 7144 6734
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 6610 7236 6666
rect 7208 6582 7328 6610
rect 7300 6254 7328 6582
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6564 4814 6684 4842
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5724 4616 5776 4622
rect 6092 4616 6144 4622
rect 5724 4558 5776 4564
rect 5828 4576 6092 4604
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4214 4660 4422
rect 4761 4380 5069 4389
rect 4761 4378 4767 4380
rect 4823 4378 4847 4380
rect 4903 4378 4927 4380
rect 4983 4378 5007 4380
rect 5063 4378 5069 4380
rect 4823 4326 4825 4378
rect 5005 4326 5007 4378
rect 4761 4324 4767 4326
rect 4823 4324 4847 4326
rect 4903 4324 4927 4326
rect 4983 4324 5007 4326
rect 5063 4324 5069 4326
rect 4761 4315 5069 4324
rect 5552 4282 5580 4558
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 4620 4208 4672 4214
rect 3698 4176 3754 4185
rect 4620 4150 4672 4156
rect 3698 4111 3754 4120
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 4101 3836 4409 3845
rect 4101 3834 4107 3836
rect 4163 3834 4187 3836
rect 4243 3834 4267 3836
rect 4323 3834 4347 3836
rect 4403 3834 4409 3836
rect 4163 3782 4165 3834
rect 4345 3782 4347 3834
rect 4101 3780 4107 3782
rect 4163 3780 4187 3782
rect 4243 3780 4267 3782
rect 4323 3780 4347 3782
rect 4403 3780 4409 3782
rect 4101 3771 4409 3780
rect 5460 3534 5488 4014
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5552 3602 5580 3946
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5644 3534 5672 4082
rect 5736 4010 5764 4558
rect 5828 4486 5856 4576
rect 6092 4558 6144 4564
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 4896 3528 4948 3534
rect 4894 3496 4896 3505
rect 5448 3528 5500 3534
rect 4948 3496 4950 3505
rect 5448 3470 5500 3476
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 4894 3431 4950 3440
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 2990 4660 3334
rect 4761 3292 5069 3301
rect 4761 3290 4767 3292
rect 4823 3290 4847 3292
rect 4903 3290 4927 3292
rect 4983 3290 5007 3292
rect 5063 3290 5069 3292
rect 4823 3238 4825 3290
rect 5005 3238 5007 3290
rect 4761 3236 4767 3238
rect 4823 3236 4847 3238
rect 4903 3236 4927 3238
rect 4983 3236 5007 3238
rect 5063 3236 5069 3238
rect 4761 3227 5069 3236
rect 5644 3126 5672 3470
rect 5828 3194 5856 4422
rect 6196 4026 6224 4762
rect 6564 4486 6592 4814
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6564 4078 6592 4422
rect 7116 4214 7144 5714
rect 7208 5370 7236 5782
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7300 5250 7328 6190
rect 7392 6186 7420 6938
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5846 7604 6054
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7668 5778 7696 6326
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7668 5658 7696 5714
rect 7852 5710 7880 6598
rect 8128 5914 8156 7346
rect 8956 6458 8984 7346
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7840 5704 7892 5710
rect 7668 5630 7788 5658
rect 7840 5646 7892 5652
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7208 5222 7328 5250
rect 7564 5228 7616 5234
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 6104 3998 6224 4026
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6368 4004 6420 4010
rect 6104 3942 6132 3998
rect 6368 3946 6420 3952
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4101 2748 4409 2757
rect 4101 2746 4107 2748
rect 4163 2746 4187 2748
rect 4243 2746 4267 2748
rect 4323 2746 4347 2748
rect 4403 2746 4409 2748
rect 4163 2694 4165 2746
rect 4345 2694 4347 2746
rect 4101 2692 4107 2694
rect 4163 2692 4187 2694
rect 4243 2692 4267 2694
rect 4323 2692 4347 2694
rect 4403 2692 4409 2694
rect 4101 2683 4409 2692
rect 6012 2650 6040 3402
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6196 2446 6224 3878
rect 6380 3126 6408 3946
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6656 2922 6684 3878
rect 6748 3194 6776 4150
rect 6828 4140 6880 4146
rect 6880 4100 7052 4128
rect 6828 4082 6880 4088
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6932 3670 6960 3946
rect 7024 3890 7052 4100
rect 7116 4078 7144 4150
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7208 3942 7236 5222
rect 7564 5170 7616 5176
rect 7576 5030 7604 5170
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7668 4622 7696 5510
rect 7760 5250 7788 5630
rect 7852 5370 7880 5646
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7760 5234 7880 5250
rect 7760 5228 7892 5234
rect 7760 5222 7840 5228
rect 7840 5170 7892 5176
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7668 4214 7696 4422
rect 7760 4282 7788 4422
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7196 3936 7248 3942
rect 7024 3884 7196 3890
rect 7024 3878 7248 3884
rect 7024 3862 7236 3878
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7208 3534 7236 3862
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7470 3496 7526 3505
rect 7668 3466 7696 4150
rect 7852 3942 7880 4762
rect 7944 4622 7972 5034
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7944 4146 7972 4558
rect 8128 4146 8156 5850
rect 8312 5778 8340 6258
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8588 5846 8616 6122
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8312 5574 8340 5714
rect 8772 5642 8800 6054
rect 8864 5778 8892 6054
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3738 7880 3878
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7944 3602 7972 4082
rect 8128 3670 8156 4082
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 8220 3466 8248 4150
rect 8404 4146 8432 4422
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8496 3942 8524 4558
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 7470 3431 7526 3440
rect 7656 3460 7708 3466
rect 7484 3398 7512 3431
rect 7656 3402 7708 3408
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 8680 3058 8708 3606
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8772 3194 8800 3402
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 9140 2650 9168 8910
rect 9508 8634 9536 9522
rect 10336 9382 10364 13874
rect 10888 13870 10916 14418
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10403 13628 10711 13637
rect 10403 13626 10409 13628
rect 10465 13626 10489 13628
rect 10545 13626 10569 13628
rect 10625 13626 10649 13628
rect 10705 13626 10711 13628
rect 10465 13574 10467 13626
rect 10647 13574 10649 13626
rect 10403 13572 10409 13574
rect 10465 13572 10489 13574
rect 10545 13572 10569 13574
rect 10625 13572 10649 13574
rect 10705 13572 10711 13574
rect 10403 13563 10711 13572
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10403 12540 10711 12549
rect 10403 12538 10409 12540
rect 10465 12538 10489 12540
rect 10545 12538 10569 12540
rect 10625 12538 10649 12540
rect 10705 12538 10711 12540
rect 10465 12486 10467 12538
rect 10647 12486 10649 12538
rect 10403 12484 10409 12486
rect 10465 12484 10489 12486
rect 10545 12484 10569 12486
rect 10625 12484 10649 12486
rect 10705 12484 10711 12486
rect 10403 12475 10711 12484
rect 10796 11898 10824 13194
rect 10888 12918 10916 13262
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10980 12434 11008 14758
rect 11348 14414 11376 14894
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11063 14172 11371 14181
rect 11063 14170 11069 14172
rect 11125 14170 11149 14172
rect 11205 14170 11229 14172
rect 11285 14170 11309 14172
rect 11365 14170 11371 14172
rect 11125 14118 11127 14170
rect 11307 14118 11309 14170
rect 11063 14116 11069 14118
rect 11125 14116 11149 14118
rect 11205 14116 11229 14118
rect 11285 14116 11309 14118
rect 11365 14116 11371 14118
rect 11063 14107 11371 14116
rect 11063 13084 11371 13093
rect 11063 13082 11069 13084
rect 11125 13082 11149 13084
rect 11205 13082 11229 13084
rect 11285 13082 11309 13084
rect 11365 13082 11371 13084
rect 11125 13030 11127 13082
rect 11307 13030 11309 13082
rect 11063 13028 11069 13030
rect 11125 13028 11149 13030
rect 11205 13028 11229 13030
rect 11285 13028 11309 13030
rect 11365 13028 11371 13030
rect 11063 13019 11371 13028
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10888 12406 11008 12434
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10403 11452 10711 11461
rect 10403 11450 10409 11452
rect 10465 11450 10489 11452
rect 10545 11450 10569 11452
rect 10625 11450 10649 11452
rect 10705 11450 10711 11452
rect 10465 11398 10467 11450
rect 10647 11398 10649 11450
rect 10403 11396 10409 11398
rect 10465 11396 10489 11398
rect 10545 11396 10569 11398
rect 10625 11396 10649 11398
rect 10705 11396 10711 11398
rect 10403 11387 10711 11396
rect 10888 10674 10916 12406
rect 11072 12152 11100 12786
rect 10980 12124 11100 12152
rect 10980 11880 11008 12124
rect 11063 11996 11371 12005
rect 11063 11994 11069 11996
rect 11125 11994 11149 11996
rect 11205 11994 11229 11996
rect 11285 11994 11309 11996
rect 11365 11994 11371 11996
rect 11125 11942 11127 11994
rect 11307 11942 11309 11994
rect 11063 11940 11069 11942
rect 11125 11940 11149 11942
rect 11205 11940 11229 11942
rect 11285 11940 11309 11942
rect 11365 11940 11371 11942
rect 11063 11931 11371 11940
rect 10980 11852 11100 11880
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10980 11150 11008 11562
rect 11072 11354 11100 11852
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10403 10364 10711 10373
rect 10403 10362 10409 10364
rect 10465 10362 10489 10364
rect 10545 10362 10569 10364
rect 10625 10362 10649 10364
rect 10705 10362 10711 10364
rect 10465 10310 10467 10362
rect 10647 10310 10649 10362
rect 10403 10308 10409 10310
rect 10465 10308 10489 10310
rect 10545 10308 10569 10310
rect 10625 10308 10649 10310
rect 10705 10308 10711 10310
rect 10403 10299 10711 10308
rect 10980 10062 11008 11086
rect 11063 10908 11371 10917
rect 11063 10906 11069 10908
rect 11125 10906 11149 10908
rect 11205 10906 11229 10908
rect 11285 10906 11309 10908
rect 11365 10906 11371 10908
rect 11125 10854 11127 10906
rect 11307 10854 11309 10906
rect 11063 10852 11069 10854
rect 11125 10852 11149 10854
rect 11205 10852 11229 10854
rect 11285 10852 11309 10854
rect 11365 10852 11371 10854
rect 11063 10843 11371 10852
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10403 9276 10711 9285
rect 10403 9274 10409 9276
rect 10465 9274 10489 9276
rect 10545 9274 10569 9276
rect 10625 9274 10649 9276
rect 10705 9274 10711 9276
rect 10465 9222 10467 9274
rect 10647 9222 10649 9274
rect 10403 9220 10409 9222
rect 10465 9220 10489 9222
rect 10545 9220 10569 9222
rect 10625 9220 10649 9222
rect 10705 9220 10711 9222
rect 10403 9211 10711 9220
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 10152 8090 10180 8842
rect 10888 8498 10916 9522
rect 10980 9518 11008 9998
rect 11063 9820 11371 9829
rect 11063 9818 11069 9820
rect 11125 9818 11149 9820
rect 11205 9818 11229 9820
rect 11285 9818 11309 9820
rect 11365 9818 11371 9820
rect 11125 9766 11127 9818
rect 11307 9766 11309 9818
rect 11063 9764 11069 9766
rect 11125 9764 11149 9766
rect 11205 9764 11229 9766
rect 11285 9764 11309 9766
rect 11365 9764 11371 9766
rect 11063 9755 11371 9764
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 11063 8732 11371 8741
rect 11063 8730 11069 8732
rect 11125 8730 11149 8732
rect 11205 8730 11229 8732
rect 11285 8730 11309 8732
rect 11365 8730 11371 8732
rect 11125 8678 11127 8730
rect 11307 8678 11309 8730
rect 11063 8676 11069 8678
rect 11125 8676 11149 8678
rect 11205 8676 11229 8678
rect 11285 8676 11309 8678
rect 11365 8676 11371 8678
rect 11063 8667 11371 8676
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10403 8188 10711 8197
rect 10403 8186 10409 8188
rect 10465 8186 10489 8188
rect 10545 8186 10569 8188
rect 10625 8186 10649 8188
rect 10705 8186 10711 8188
rect 10465 8134 10467 8186
rect 10647 8134 10649 8186
rect 10403 8132 10409 8134
rect 10465 8132 10489 8134
rect 10545 8132 10569 8134
rect 10625 8132 10649 8134
rect 10705 8132 10711 8134
rect 10403 8123 10711 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 7206 9260 7822
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9232 6458 9260 7142
rect 9600 6866 9628 7142
rect 9784 7002 9812 7210
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9324 6458 9352 6666
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9232 4078 9260 6394
rect 9324 6322 9352 6394
rect 9416 6322 9444 6598
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9692 6186 9720 6598
rect 9876 6458 9904 7686
rect 10060 7546 10088 7754
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10152 7478 10180 7890
rect 10244 7546 10272 7958
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10152 6458 10180 7414
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10244 6458 10272 7278
rect 10336 6866 10364 7686
rect 10403 7100 10711 7109
rect 10403 7098 10409 7100
rect 10465 7098 10489 7100
rect 10545 7098 10569 7100
rect 10625 7098 10649 7100
rect 10705 7098 10711 7100
rect 10465 7046 10467 7098
rect 10647 7046 10649 7098
rect 10403 7044 10409 7046
rect 10465 7044 10489 7046
rect 10545 7044 10569 7046
rect 10625 7044 10649 7046
rect 10705 7044 10711 7046
rect 10403 7035 10711 7044
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9588 5840 9640 5846
rect 9640 5788 9812 5794
rect 9588 5782 9812 5788
rect 9600 5766 9812 5782
rect 9784 5710 9812 5766
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9508 4282 9536 5102
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9876 4146 9904 6394
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9968 5914 9996 6258
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10060 5914 10088 6122
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10244 5710 10272 6258
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10336 5710 10364 6190
rect 10403 6012 10711 6021
rect 10403 6010 10409 6012
rect 10465 6010 10489 6012
rect 10545 6010 10569 6012
rect 10625 6010 10649 6012
rect 10705 6010 10711 6012
rect 10465 5958 10467 6010
rect 10647 5958 10649 6010
rect 10403 5956 10409 5958
rect 10465 5956 10489 5958
rect 10545 5956 10569 5958
rect 10625 5956 10649 5958
rect 10705 5956 10711 5958
rect 10403 5947 10711 5956
rect 10796 5846 10824 6190
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10336 5234 10364 5646
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10796 5166 10824 5646
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10403 4924 10711 4933
rect 10403 4922 10409 4924
rect 10465 4922 10489 4924
rect 10545 4922 10569 4924
rect 10625 4922 10649 4924
rect 10705 4922 10711 4924
rect 10465 4870 10467 4922
rect 10647 4870 10649 4922
rect 10403 4868 10409 4870
rect 10465 4868 10489 4870
rect 10545 4868 10569 4870
rect 10625 4868 10649 4870
rect 10705 4868 10711 4870
rect 10403 4859 10711 4868
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10060 4214 10088 4490
rect 10796 4214 10824 5102
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9232 3738 9260 4014
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9968 3058 9996 3470
rect 10060 3126 10088 3878
rect 10403 3836 10711 3845
rect 10403 3834 10409 3836
rect 10465 3834 10489 3836
rect 10545 3834 10569 3836
rect 10625 3834 10649 3836
rect 10705 3834 10711 3836
rect 10465 3782 10467 3834
rect 10647 3782 10649 3834
rect 10403 3780 10409 3782
rect 10465 3780 10489 3782
rect 10545 3780 10569 3782
rect 10625 3780 10649 3782
rect 10705 3780 10711 3782
rect 10403 3771 10711 3780
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10403 2748 10711 2757
rect 10403 2746 10409 2748
rect 10465 2746 10489 2748
rect 10545 2746 10569 2748
rect 10625 2746 10649 2748
rect 10705 2746 10711 2748
rect 10465 2694 10467 2746
rect 10647 2694 10649 2746
rect 10403 2692 10409 2694
rect 10465 2692 10489 2694
rect 10545 2692 10569 2694
rect 10625 2692 10649 2694
rect 10705 2692 10711 2694
rect 10403 2683 10711 2692
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 3896 800 3924 2382
rect 4761 2204 5069 2213
rect 4761 2202 4767 2204
rect 4823 2202 4847 2204
rect 4903 2202 4927 2204
rect 4983 2202 5007 2204
rect 5063 2202 5069 2204
rect 4823 2150 4825 2202
rect 5005 2150 5007 2202
rect 4761 2148 4767 2150
rect 4823 2148 4847 2150
rect 4903 2148 4927 2150
rect 4983 2148 5007 2150
rect 5063 2148 5069 2150
rect 4761 2139 5069 2148
rect 7760 800 7788 2382
rect 10888 2310 10916 8434
rect 11063 7644 11371 7653
rect 11063 7642 11069 7644
rect 11125 7642 11149 7644
rect 11205 7642 11229 7644
rect 11285 7642 11309 7644
rect 11365 7642 11371 7644
rect 11125 7590 11127 7642
rect 11307 7590 11309 7642
rect 11063 7588 11069 7590
rect 11125 7588 11149 7590
rect 11205 7588 11229 7590
rect 11285 7588 11309 7590
rect 11365 7588 11371 7590
rect 11063 7579 11371 7588
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 7018 11192 7142
rect 10980 7002 11192 7018
rect 10968 6996 11192 7002
rect 11020 6990 11192 6996
rect 10968 6938 11020 6944
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10980 6322 11008 6666
rect 11063 6556 11371 6565
rect 11063 6554 11069 6556
rect 11125 6554 11149 6556
rect 11205 6554 11229 6556
rect 11285 6554 11309 6556
rect 11365 6554 11371 6556
rect 11125 6502 11127 6554
rect 11307 6502 11309 6554
rect 11063 6500 11069 6502
rect 11125 6500 11149 6502
rect 11205 6500 11229 6502
rect 11285 6500 11309 6502
rect 11365 6500 11371 6502
rect 11063 6491 11371 6500
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11072 5914 11100 6190
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11348 5846 11376 6054
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 10980 5630 11100 5658
rect 10980 5250 11008 5630
rect 11072 5574 11100 5630
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11063 5468 11371 5477
rect 11063 5466 11069 5468
rect 11125 5466 11149 5468
rect 11205 5466 11229 5468
rect 11285 5466 11309 5468
rect 11365 5466 11371 5468
rect 11125 5414 11127 5466
rect 11307 5414 11309 5466
rect 11063 5412 11069 5414
rect 11125 5412 11149 5414
rect 11205 5412 11229 5414
rect 11285 5412 11309 5414
rect 11365 5412 11371 5414
rect 11063 5403 11371 5412
rect 10980 5222 11192 5250
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10980 4826 11008 4966
rect 11072 4826 11100 5102
rect 11164 5030 11192 5222
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10980 4486 11008 4762
rect 11060 4616 11112 4622
rect 11164 4604 11192 4966
rect 11112 4576 11192 4604
rect 11060 4558 11112 4564
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10980 4146 11008 4422
rect 11063 4380 11371 4389
rect 11063 4378 11069 4380
rect 11125 4378 11149 4380
rect 11205 4378 11229 4380
rect 11285 4378 11309 4380
rect 11365 4378 11371 4380
rect 11125 4326 11127 4378
rect 11307 4326 11309 4378
rect 11063 4324 11069 4326
rect 11125 4324 11149 4326
rect 11205 4324 11229 4326
rect 11285 4324 11309 4326
rect 11365 4324 11371 4326
rect 11063 4315 11371 4324
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 4010 11192 4082
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 3534 11100 3878
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11063 3292 11371 3301
rect 11063 3290 11069 3292
rect 11125 3290 11149 3292
rect 11205 3290 11229 3292
rect 11285 3290 11309 3292
rect 11365 3290 11371 3292
rect 11125 3238 11127 3290
rect 11307 3238 11309 3290
rect 11063 3236 11069 3238
rect 11125 3236 11149 3238
rect 11205 3236 11229 3238
rect 11285 3236 11309 3238
rect 11365 3236 11371 3238
rect 11063 3227 11371 3236
rect 11440 2514 11468 16476
rect 11532 16250 11560 16526
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11532 14074 11560 14214
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13274 11560 13670
rect 11624 13394 11652 14418
rect 11716 13954 11744 18022
rect 11808 17610 11836 18158
rect 11900 17814 11928 18226
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11808 17134 11836 17546
rect 11900 17134 11928 17750
rect 12084 17746 12112 19382
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 12084 16726 12112 17682
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 12084 16454 12112 16662
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11900 15162 11928 15438
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 12084 14958 12112 16390
rect 12176 15162 12204 19246
rect 12452 17678 12480 20470
rect 13280 20330 13308 20878
rect 14278 20839 14334 20848
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 12636 19174 12664 19926
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12728 19514 12756 19790
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18290 12664 19110
rect 12728 18698 12756 19450
rect 12820 19446 12848 19654
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 13280 18766 13308 20266
rect 13464 19854 13492 20402
rect 13648 19922 13676 20402
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13648 19446 13676 19858
rect 14004 19780 14056 19786
rect 14004 19722 14056 19728
rect 14016 19514 14044 19722
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12912 17610 12940 18566
rect 13004 18086 13032 18702
rect 13648 18698 13676 19382
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13648 18578 13676 18634
rect 13556 18550 13676 18578
rect 13556 18290 13584 18550
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 13096 17898 13124 18090
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13096 17882 13216 17898
rect 13096 17876 13228 17882
rect 13096 17870 13176 17876
rect 13176 17818 13228 17824
rect 13372 17610 13400 18022
rect 13832 17814 13860 18022
rect 13924 17882 13952 18226
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13728 17672 13780 17678
rect 14108 17626 14136 19654
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18970 14320 19110
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 13728 17614 13780 17620
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12452 15706 12480 16458
rect 12544 16114 12572 17478
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16250 12756 17070
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12624 15088 12676 15094
rect 12622 15056 12624 15065
rect 12676 15056 12678 15065
rect 12532 15020 12584 15026
rect 12622 14991 12678 15000
rect 12532 14962 12584 14968
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11808 14074 11836 14894
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11900 14006 11928 14486
rect 12084 14482 12112 14894
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12268 14074 12296 14758
rect 12452 14482 12480 14758
rect 12544 14618 12572 14962
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 11888 14000 11940 14006
rect 11716 13926 11836 13954
rect 11888 13942 11940 13948
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11716 13308 11744 13738
rect 11808 13734 11836 13926
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11796 13320 11848 13326
rect 11716 13280 11796 13308
rect 11532 13246 11652 13274
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11532 12850 11560 13126
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11624 12646 11652 13246
rect 11716 12782 11744 13280
rect 11796 13262 11848 13268
rect 11900 12850 11928 13806
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11532 11898 11560 12242
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 10062 11560 11494
rect 11624 11354 11652 12174
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11716 11218 11744 12718
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 11778 11836 12582
rect 11900 12238 11928 12786
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11808 11750 11928 11778
rect 11992 11762 12020 14010
rect 12360 13326 12388 14282
rect 12636 13530 12664 14826
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12084 11762 12112 13194
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12176 12442 12204 12718
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11354 11836 11630
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11900 11150 11928 11750
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12176 11354 12204 11562
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11716 10810 11744 11018
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9178 11560 9998
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11716 8974 11744 9590
rect 11900 9178 11928 11086
rect 11992 10266 12020 11222
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12164 9580 12216 9586
rect 12084 9540 12164 9568
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 5574 11560 7142
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 4758 11560 5510
rect 11624 5370 11652 6190
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11532 4214 11560 4694
rect 11624 4214 11652 4966
rect 11716 4758 11744 8910
rect 11900 8294 11928 9114
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8566 12020 8774
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 12084 8498 12112 9540
rect 12164 9522 12216 9528
rect 12360 9382 12388 13262
rect 12728 12434 12756 15982
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12820 14074 12848 14418
rect 12912 14074 12940 17546
rect 13372 15858 13400 17546
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 16250 13492 16594
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13372 15830 13492 15858
rect 13464 14278 13492 15830
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13464 13394 13492 14214
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12986 12848 13262
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12912 12918 12940 13126
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12728 12406 13032 12434
rect 13004 11694 13032 12406
rect 13096 11762 13124 12922
rect 13556 12442 13584 17546
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13648 16726 13676 17002
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13648 15366 13676 16662
rect 13740 15638 13768 17614
rect 13832 17598 14136 17626
rect 14200 17610 14228 18634
rect 14292 17882 14320 18906
rect 14464 18896 14516 18902
rect 14462 18864 14464 18873
rect 14516 18864 14518 18873
rect 14462 18799 14518 18808
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14188 17604 14240 17610
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13740 15162 13768 15574
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13648 13326 13676 13874
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13188 11898 13216 12106
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12452 9654 12480 11086
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 10130 12848 10474
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12544 9586 12572 9998
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12636 9058 12664 9998
rect 12808 9988 12860 9994
rect 12452 9042 12664 9058
rect 12440 9036 12664 9042
rect 12492 9030 12664 9036
rect 12440 8978 12492 8984
rect 12636 8974 12664 9030
rect 12728 9948 12808 9976
rect 12256 8968 12308 8974
rect 12624 8968 12676 8974
rect 12308 8916 12480 8922
rect 12256 8910 12480 8916
rect 12624 8910 12676 8916
rect 12268 8894 12480 8910
rect 12452 8566 12480 8894
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11808 7546 11836 7754
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11900 6662 11928 7346
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6458 12020 6598
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 4282 11928 4626
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11624 3194 11652 4150
rect 11992 4146 12020 5510
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11992 3738 12020 4082
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 12084 2650 12112 8434
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 7478 12296 8230
rect 12452 7886 12480 8298
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12268 7002 12296 7414
rect 12728 7410 12756 9948
rect 12808 9930 12860 9936
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12820 9178 12848 9454
rect 12912 9450 12940 9522
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8566 12848 8978
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12912 8090 12940 9386
rect 13004 9178 13032 11630
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10674 13676 10950
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 13096 9042 13124 10474
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 10062 13216 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13372 10130 13492 10146
rect 13360 10124 13492 10130
rect 13412 10118 13492 10124
rect 13360 10066 13412 10072
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 9654 13216 9862
rect 13372 9722 13400 9930
rect 13464 9874 13492 10118
rect 13556 10062 13584 10202
rect 13648 10062 13676 10610
rect 13740 10198 13768 15098
rect 13832 11150 13860 17598
rect 14188 17546 14240 17552
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13924 14618 13952 17478
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 14016 16794 14044 17206
rect 14200 17134 14228 17546
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14188 16992 14240 16998
rect 14292 16946 14320 17818
rect 14240 16940 14320 16946
rect 14188 16934 14320 16940
rect 14200 16918 14320 16934
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14384 16658 14412 18702
rect 14568 18426 14596 18906
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14646 18320 14702 18329
rect 14646 18255 14648 18264
rect 14700 18255 14702 18264
rect 14648 18226 14700 18232
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14568 17202 14596 18022
rect 14752 17626 14780 21490
rect 15212 21434 15240 22442
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 15304 21554 15332 21966
rect 15580 21554 15608 22374
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15120 21418 15240 21434
rect 15108 21412 15240 21418
rect 15160 21406 15240 21412
rect 15108 21354 15160 21360
rect 15212 21010 15240 21406
rect 15580 21350 15608 21490
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15856 20874 15884 25706
rect 16304 25696 16356 25702
rect 16304 25638 16356 25644
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 16040 24410 16068 25230
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 16316 24256 16344 25638
rect 16396 25356 16448 25362
rect 16396 25298 16448 25304
rect 16408 24750 16436 25298
rect 16592 24954 16620 26318
rect 17420 26246 17448 26318
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17408 26240 17460 26246
rect 17408 26182 17460 26188
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 16705 25596 17013 25605
rect 16705 25594 16711 25596
rect 16767 25594 16791 25596
rect 16847 25594 16871 25596
rect 16927 25594 16951 25596
rect 17007 25594 17013 25596
rect 16767 25542 16769 25594
rect 16949 25542 16951 25594
rect 16705 25540 16711 25542
rect 16767 25540 16791 25542
rect 16847 25540 16871 25542
rect 16927 25540 16951 25542
rect 17007 25540 17013 25542
rect 16705 25531 17013 25540
rect 17052 25362 17080 25774
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16776 24818 16804 25094
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16408 24410 16436 24550
rect 16396 24404 16448 24410
rect 16396 24346 16448 24352
rect 16500 24290 16528 24686
rect 16592 24410 16620 24754
rect 16960 24698 16988 25230
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24818 17080 25094
rect 17144 24954 17172 25842
rect 17236 25294 17264 26182
rect 17365 26140 17673 26149
rect 17365 26138 17371 26140
rect 17427 26138 17451 26140
rect 17507 26138 17531 26140
rect 17587 26138 17611 26140
rect 17667 26138 17673 26140
rect 17427 26086 17429 26138
rect 17609 26086 17611 26138
rect 17365 26084 17371 26086
rect 17427 26084 17451 26086
rect 17507 26084 17531 26086
rect 17587 26084 17611 26086
rect 17667 26084 17673 26086
rect 17365 26075 17673 26084
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17236 24954 17264 25094
rect 17365 25052 17673 25061
rect 17365 25050 17371 25052
rect 17427 25050 17451 25052
rect 17507 25050 17531 25052
rect 17587 25050 17611 25052
rect 17667 25050 17673 25052
rect 17427 24998 17429 25050
rect 17609 24998 17611 25050
rect 17365 24996 17371 24998
rect 17427 24996 17451 24998
rect 17507 24996 17531 24998
rect 17587 24996 17611 24998
rect 17667 24996 17673 24998
rect 17365 24987 17673 24996
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17788 24857 17816 26318
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17130 24848 17186 24857
rect 17040 24812 17092 24818
rect 17774 24848 17830 24857
rect 17130 24783 17132 24792
rect 17040 24754 17092 24760
rect 17184 24783 17186 24792
rect 17224 24812 17276 24818
rect 17132 24754 17184 24760
rect 17224 24754 17276 24760
rect 17316 24812 17368 24818
rect 17774 24783 17830 24792
rect 17316 24754 17368 24760
rect 16960 24670 17080 24698
rect 16705 24508 17013 24517
rect 16705 24506 16711 24508
rect 16767 24506 16791 24508
rect 16847 24506 16871 24508
rect 16927 24506 16951 24508
rect 17007 24506 17013 24508
rect 16767 24454 16769 24506
rect 16949 24454 16951 24506
rect 16705 24452 16711 24454
rect 16767 24452 16791 24454
rect 16847 24452 16871 24454
rect 16927 24452 16951 24454
rect 17007 24452 17013 24454
rect 16705 24443 17013 24452
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 17052 24342 17080 24670
rect 17236 24342 17264 24754
rect 17328 24614 17356 24754
rect 17880 24682 17908 25434
rect 18248 24818 18276 25638
rect 18432 24818 18460 26386
rect 19064 26376 19116 26382
rect 19064 26318 19116 26324
rect 18788 26240 18840 26246
rect 18788 26182 18840 26188
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18708 24818 18736 25978
rect 18800 25702 18828 26182
rect 19076 25838 19104 26318
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18800 24886 18828 25638
rect 18880 25152 18932 25158
rect 18880 25094 18932 25100
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 18892 24818 18920 25094
rect 19076 24818 19104 25774
rect 19156 25220 19208 25226
rect 19156 25162 19208 25168
rect 19168 24818 19196 25162
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 17500 24676 17552 24682
rect 17500 24618 17552 24624
rect 17868 24676 17920 24682
rect 17868 24618 17920 24624
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17040 24336 17092 24342
rect 16396 24268 16448 24274
rect 16316 24228 16396 24256
rect 16316 23798 16344 24228
rect 16500 24262 16620 24290
rect 17040 24278 17092 24284
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 16396 24210 16448 24216
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15948 22234 15976 22986
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16028 22500 16080 22506
rect 16028 22442 16080 22448
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 16040 21962 16068 22442
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16132 22098 16160 22374
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16224 22030 16252 22918
rect 16316 22710 16344 23734
rect 16500 23526 16528 24142
rect 16592 23866 16620 24262
rect 17052 24206 17080 24278
rect 17512 24274 17540 24618
rect 17972 24410 18000 24754
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 17365 23964 17673 23973
rect 17365 23962 17371 23964
rect 17427 23962 17451 23964
rect 17507 23962 17531 23964
rect 17587 23962 17611 23964
rect 17667 23962 17673 23964
rect 17427 23910 17429 23962
rect 17609 23910 17611 23962
rect 17365 23908 17371 23910
rect 17427 23908 17451 23910
rect 17507 23908 17531 23910
rect 17587 23908 17611 23910
rect 17667 23908 17673 23910
rect 17365 23899 17673 23908
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 16705 23420 17013 23429
rect 16705 23418 16711 23420
rect 16767 23418 16791 23420
rect 16847 23418 16871 23420
rect 16927 23418 16951 23420
rect 17007 23418 17013 23420
rect 16767 23366 16769 23418
rect 16949 23366 16951 23418
rect 16705 23364 16711 23366
rect 16767 23364 16791 23366
rect 16847 23364 16871 23366
rect 16927 23364 16951 23366
rect 17007 23364 17013 23366
rect 16705 23355 17013 23364
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16304 22704 16356 22710
rect 16304 22646 16356 22652
rect 16408 22642 16436 23054
rect 17052 22710 17080 23462
rect 17972 23186 18000 24346
rect 18156 24206 18184 24754
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18052 23248 18104 23254
rect 18052 23190 18104 23196
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16408 22522 16436 22578
rect 17144 22574 17172 22918
rect 17365 22876 17673 22885
rect 17365 22874 17371 22876
rect 17427 22874 17451 22876
rect 17507 22874 17531 22876
rect 17587 22874 17611 22876
rect 17667 22874 17673 22876
rect 17427 22822 17429 22874
rect 17609 22822 17611 22874
rect 17365 22820 17371 22822
rect 17427 22820 17451 22822
rect 17507 22820 17531 22822
rect 17587 22820 17611 22822
rect 17667 22820 17673 22822
rect 17365 22811 17673 22820
rect 16316 22494 16436 22522
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 16316 22438 16344 22494
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15198 20496 15254 20505
rect 15198 20431 15200 20440
rect 15252 20431 15254 20440
rect 15200 20402 15252 20408
rect 16040 20262 16068 21286
rect 16132 21010 16160 21558
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 14832 18692 14884 18698
rect 14832 18634 14884 18640
rect 14844 18290 14872 18634
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 14752 17598 14872 17626
rect 14844 17542 14872 17598
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14752 17338 14780 17478
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14384 14414 14412 16594
rect 14660 16046 14688 16934
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14476 14618 14504 15438
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 11762 14136 13262
rect 14292 12986 14320 14282
rect 14384 13938 14412 14350
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13924 10130 13952 10406
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 14384 10062 14412 10610
rect 14476 10062 14504 13806
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11830 14596 12038
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13464 9846 13676 9874
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13188 9382 13216 9590
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13280 9178 13308 9522
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8498 13124 8842
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13188 8106 13216 9114
rect 13648 9110 13676 9846
rect 13832 9450 13860 9930
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 14108 9178 14136 9522
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13452 9104 13504 9110
rect 13636 9104 13688 9110
rect 13504 9052 13636 9058
rect 13452 9046 13688 9052
rect 13268 9036 13320 9042
rect 13464 9030 13676 9046
rect 13268 8978 13320 8984
rect 13280 8294 13308 8978
rect 14016 8974 14044 9114
rect 14200 9110 14228 9386
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8498 13400 8774
rect 13464 8634 13492 8842
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13464 8498 13492 8570
rect 14384 8566 14412 9522
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 12900 8084 12952 8090
rect 13188 8078 13400 8106
rect 13924 8090 13952 8434
rect 14568 8294 14596 9862
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 12900 8026 12952 8032
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12176 6458 12204 6666
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12268 6390 12296 6938
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12452 6322 12480 7346
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 6390 12756 6734
rect 12912 6730 12940 6802
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12912 6322 12940 6666
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12636 4146 12664 4558
rect 12820 4146 12848 5714
rect 12912 5710 12940 6258
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12452 3534 12480 3674
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 12820 2446 12848 4082
rect 12912 3602 12940 5646
rect 13188 5642 13216 6598
rect 13280 6322 13308 6598
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12912 2990 12940 3538
rect 13004 3466 13032 3878
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13096 3058 13124 3334
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 13372 2774 13400 8078
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14200 5914 14228 6326
rect 14384 6118 14412 6734
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 13728 4616 13780 4622
rect 13912 4616 13964 4622
rect 13728 4558 13780 4564
rect 13910 4584 13912 4593
rect 13964 4584 13966 4593
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13648 4282 13676 4490
rect 13740 4282 13768 4558
rect 13910 4519 13966 4528
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13648 3466 13676 4218
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 14016 3398 14044 4490
rect 14108 4146 14136 5782
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 3534 14136 4082
rect 14200 4078 14228 4966
rect 14292 4146 14320 5170
rect 14384 5166 14412 6054
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14384 4214 14412 5102
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14476 4282 14504 4558
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14292 3670 14320 4082
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14280 3664 14332 3670
rect 14280 3606 14332 3612
rect 14384 3602 14412 3878
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14568 3534 14596 4694
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13372 2746 13492 2774
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 11063 2204 11371 2213
rect 11063 2202 11069 2204
rect 11125 2202 11149 2204
rect 11205 2202 11229 2204
rect 11285 2202 11309 2204
rect 11365 2202 11371 2204
rect 11125 2150 11127 2202
rect 11307 2150 11309 2202
rect 11063 2148 11069 2150
rect 11125 2148 11149 2150
rect 11205 2148 11229 2150
rect 11285 2148 11309 2150
rect 11365 2148 11371 2150
rect 11063 2139 11371 2148
rect 11624 800 11652 2382
rect 13464 2378 13492 2746
rect 13832 2650 13860 3062
rect 14660 2774 14688 15982
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 14346 14780 14894
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10266 14780 10950
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14844 9042 14872 11834
rect 15028 11150 15056 18022
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16182 15148 16934
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10674 14964 10950
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14936 9586 14964 9998
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 15120 9081 15148 16118
rect 15212 14550 15240 19450
rect 15948 19378 15976 20198
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15764 18630 15792 19246
rect 16132 18766 16160 19654
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15948 18426 15976 18702
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 16132 18193 16160 18294
rect 16118 18184 16174 18193
rect 16118 18119 16174 18128
rect 16132 17746 16160 18119
rect 16224 18086 16252 21830
rect 16316 21690 16344 22374
rect 16705 22332 17013 22341
rect 16705 22330 16711 22332
rect 16767 22330 16791 22332
rect 16847 22330 16871 22332
rect 16927 22330 16951 22332
rect 17007 22330 17013 22332
rect 16767 22278 16769 22330
rect 16949 22278 16951 22330
rect 16705 22276 16711 22278
rect 16767 22276 16791 22278
rect 16847 22276 16871 22278
rect 16927 22276 16951 22278
rect 17007 22276 17013 22278
rect 16705 22267 17013 22276
rect 17052 22094 17080 22374
rect 17236 22234 17264 22374
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 16868 22066 17080 22094
rect 16868 22030 16896 22066
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16592 20942 16620 21830
rect 16868 21486 16896 21966
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16705 21244 17013 21253
rect 16705 21242 16711 21244
rect 16767 21242 16791 21244
rect 16847 21242 16871 21244
rect 16927 21242 16951 21244
rect 17007 21242 17013 21244
rect 16767 21190 16769 21242
rect 16949 21190 16951 21242
rect 16705 21188 16711 21190
rect 16767 21188 16791 21190
rect 16847 21188 16871 21190
rect 16927 21188 16951 21190
rect 17007 21188 17013 21190
rect 16705 21179 17013 21188
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 20346 16620 20742
rect 16868 20466 16896 20946
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16500 20318 16620 20346
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16316 19854 16344 20198
rect 16500 19990 16528 20318
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16592 19990 16620 20198
rect 16705 20156 17013 20165
rect 16705 20154 16711 20156
rect 16767 20154 16791 20156
rect 16847 20154 16871 20156
rect 16927 20154 16951 20156
rect 17007 20154 17013 20156
rect 16767 20102 16769 20154
rect 16949 20102 16951 20154
rect 16705 20100 16711 20102
rect 16767 20100 16791 20102
rect 16847 20100 16871 20102
rect 16927 20100 16951 20102
rect 17007 20100 17013 20102
rect 16705 20091 17013 20100
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16500 19854 16528 19926
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19242 16620 19654
rect 17052 19258 17080 21830
rect 17144 21690 17172 22170
rect 17328 22098 17356 22510
rect 17776 22500 17828 22506
rect 17776 22442 17828 22448
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17696 21842 17724 22374
rect 17788 22166 17816 22442
rect 17880 22234 17908 22986
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17776 22160 17828 22166
rect 17776 22102 17828 22108
rect 17788 22030 17816 22102
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17880 21962 17908 22170
rect 18064 22094 18092 23190
rect 18156 22778 18184 24142
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 18064 22066 18184 22094
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 18052 21956 18104 21962
rect 18052 21898 18104 21904
rect 17696 21814 17816 21842
rect 17365 21788 17673 21797
rect 17365 21786 17371 21788
rect 17427 21786 17451 21788
rect 17507 21786 17531 21788
rect 17587 21786 17611 21788
rect 17667 21786 17673 21788
rect 17427 21734 17429 21786
rect 17609 21734 17611 21786
rect 17365 21732 17371 21734
rect 17427 21732 17451 21734
rect 17507 21732 17531 21734
rect 17587 21732 17611 21734
rect 17667 21732 17673 21734
rect 17365 21723 17673 21732
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17144 20466 17172 20810
rect 17236 20534 17264 21082
rect 17512 20942 17540 21422
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17365 20700 17673 20709
rect 17365 20698 17371 20700
rect 17427 20698 17451 20700
rect 17507 20698 17531 20700
rect 17587 20698 17611 20700
rect 17667 20698 17673 20700
rect 17427 20646 17429 20698
rect 17609 20646 17611 20698
rect 17365 20644 17371 20646
rect 17427 20644 17451 20646
rect 17507 20644 17531 20646
rect 17587 20644 17611 20646
rect 17667 20644 17673 20646
rect 17365 20635 17673 20644
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17130 19816 17186 19825
rect 17130 19751 17186 19760
rect 17144 19378 17172 19751
rect 17236 19496 17264 20470
rect 17788 20398 17816 21814
rect 18064 21622 18092 21898
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17880 19854 17908 21286
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17972 20466 18000 21082
rect 18064 20942 18092 21558
rect 18156 21418 18184 22066
rect 18248 21554 18276 22918
rect 18340 22642 18368 22918
rect 18524 22642 18552 23054
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18328 22500 18380 22506
rect 18328 22442 18380 22448
rect 18340 22166 18368 22442
rect 18524 22234 18552 22578
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18328 22160 18380 22166
rect 18328 22102 18380 22108
rect 18616 21962 18644 22646
rect 18892 22438 18920 24142
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18984 21622 19012 21830
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18616 21146 18644 21490
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18052 20936 18104 20942
rect 19076 20913 19104 24754
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 19260 22642 19288 22986
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19260 22234 19288 22578
rect 19248 22228 19300 22234
rect 19248 22170 19300 22176
rect 19260 22030 19288 22170
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 18052 20878 18104 20884
rect 19062 20904 19118 20913
rect 19062 20839 19118 20848
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17365 19612 17673 19621
rect 17365 19610 17371 19612
rect 17427 19610 17451 19612
rect 17507 19610 17531 19612
rect 17587 19610 17611 19612
rect 17667 19610 17673 19612
rect 17427 19558 17429 19610
rect 17609 19558 17611 19610
rect 17365 19556 17371 19558
rect 17427 19556 17451 19558
rect 17507 19556 17531 19558
rect 17587 19556 17611 19558
rect 17667 19556 17673 19558
rect 17365 19547 17673 19556
rect 17236 19468 17448 19496
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17224 19304 17276 19310
rect 16580 19236 16632 19242
rect 17052 19230 17172 19258
rect 17224 19246 17276 19252
rect 16580 19178 16632 19184
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16705 19068 17013 19077
rect 16705 19066 16711 19068
rect 16767 19066 16791 19068
rect 16847 19066 16871 19068
rect 16927 19066 16951 19068
rect 17007 19066 17013 19068
rect 16767 19014 16769 19066
rect 16949 19014 16951 19066
rect 16705 19012 16711 19014
rect 16767 19012 16791 19014
rect 16847 19012 16871 19014
rect 16927 19012 16951 19014
rect 17007 19012 17013 19014
rect 16705 19003 17013 19012
rect 17052 18902 17080 19110
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16408 18465 16436 18634
rect 16394 18456 16450 18465
rect 16394 18391 16450 18400
rect 16500 18154 16528 18838
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16868 18290 16896 18566
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16960 18086 16988 18362
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16705 17980 17013 17989
rect 16705 17978 16711 17980
rect 16767 17978 16791 17980
rect 16847 17978 16871 17980
rect 16927 17978 16951 17980
rect 17007 17978 17013 17980
rect 16767 17926 16769 17978
rect 16949 17926 16951 17978
rect 16705 17924 16711 17926
rect 16767 17924 16791 17926
rect 16847 17924 16871 17926
rect 16927 17924 16951 17926
rect 17007 17924 17013 17926
rect 16705 17915 17013 17924
rect 17052 17882 17080 18566
rect 17144 18034 17172 19230
rect 17236 19174 17264 19246
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17236 18630 17264 19110
rect 17328 18766 17356 19178
rect 17420 19174 17448 19468
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17788 18766 17816 19654
rect 17880 19446 17908 19790
rect 17972 19446 18000 20402
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17972 18766 18000 19382
rect 18064 19378 18092 20198
rect 18248 19854 18276 20266
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18156 19242 18184 19314
rect 18248 19242 18276 19790
rect 18524 19310 18552 20198
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 17365 18524 17673 18533
rect 17365 18522 17371 18524
rect 17427 18522 17451 18524
rect 17507 18522 17531 18524
rect 17587 18522 17611 18524
rect 17667 18522 17673 18524
rect 17427 18470 17429 18522
rect 17609 18470 17611 18522
rect 17365 18468 17371 18470
rect 17427 18468 17451 18470
rect 17507 18468 17531 18470
rect 17587 18468 17611 18470
rect 17667 18468 17673 18470
rect 17222 18456 17278 18465
rect 17365 18459 17673 18468
rect 17222 18391 17278 18400
rect 17236 18154 17264 18391
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17420 18193 17448 18226
rect 17406 18184 17462 18193
rect 17224 18148 17276 18154
rect 17406 18119 17462 18128
rect 17224 18090 17276 18096
rect 17408 18080 17460 18086
rect 17144 18028 17408 18034
rect 17144 18022 17460 18028
rect 17144 18006 17448 18022
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 17144 17678 17172 18006
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17365 17436 17673 17445
rect 17365 17434 17371 17436
rect 17427 17434 17451 17436
rect 17507 17434 17531 17436
rect 17587 17434 17611 17436
rect 17667 17434 17673 17436
rect 17427 17382 17429 17434
rect 17609 17382 17611 17434
rect 17365 17380 17371 17382
rect 17427 17380 17451 17382
rect 17507 17380 17531 17382
rect 17587 17380 17611 17382
rect 17667 17380 17673 17382
rect 17365 17371 17673 17380
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15212 13190 15240 14214
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15396 12986 15424 13194
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15488 11082 15516 15506
rect 15580 15502 15608 16526
rect 16592 16114 16620 17070
rect 16705 16892 17013 16901
rect 16705 16890 16711 16892
rect 16767 16890 16791 16892
rect 16847 16890 16871 16892
rect 16927 16890 16951 16892
rect 17007 16890 17013 16892
rect 16767 16838 16769 16890
rect 16949 16838 16951 16890
rect 16705 16836 16711 16838
rect 16767 16836 16791 16838
rect 16847 16836 16871 16838
rect 16927 16836 16951 16838
rect 17007 16836 17013 16838
rect 16705 16827 17013 16836
rect 17365 16348 17673 16357
rect 17365 16346 17371 16348
rect 17427 16346 17451 16348
rect 17507 16346 17531 16348
rect 17587 16346 17611 16348
rect 17667 16346 17673 16348
rect 17427 16294 17429 16346
rect 17609 16294 17611 16346
rect 17365 16292 17371 16294
rect 17427 16292 17451 16294
rect 17507 16292 17531 16294
rect 17587 16292 17611 16294
rect 17667 16292 17673 16294
rect 17365 16283 17673 16292
rect 17788 16130 17816 18566
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 17972 17746 18000 18362
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18156 17814 18184 18294
rect 18248 18290 18276 18566
rect 18708 18426 18736 18566
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16590 18000 17206
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 17696 16102 17816 16130
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16705 15804 17013 15813
rect 16705 15802 16711 15804
rect 16767 15802 16791 15804
rect 16847 15802 16871 15804
rect 16927 15802 16951 15804
rect 17007 15802 17013 15804
rect 16767 15750 16769 15802
rect 16949 15750 16951 15802
rect 16705 15748 16711 15750
rect 16767 15748 16791 15750
rect 16847 15748 16871 15750
rect 16927 15748 16951 15750
rect 17007 15748 17013 15750
rect 16705 15739 17013 15748
rect 17052 15570 17080 15846
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15580 12850 15608 15438
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15094 15792 15302
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15948 14346 15976 15506
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 16212 14340 16264 14346
rect 16316 14328 16344 14554
rect 16264 14300 16344 14328
rect 16212 14282 16264 14288
rect 15764 13870 15792 14282
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15948 13530 15976 14282
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16316 13462 16344 13806
rect 16500 13734 16528 15438
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 15162 16896 15302
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16960 14906 16988 15506
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 17052 15162 17080 15370
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17144 15094 17172 15506
rect 17604 15502 17632 15642
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 16960 14878 17080 14906
rect 16705 14716 17013 14725
rect 16705 14714 16711 14716
rect 16767 14714 16791 14716
rect 16847 14714 16871 14716
rect 16927 14714 16951 14716
rect 17007 14714 17013 14716
rect 16767 14662 16769 14714
rect 16949 14662 16951 14714
rect 16705 14660 16711 14662
rect 16767 14660 16791 14662
rect 16847 14660 16871 14662
rect 16927 14660 16951 14662
rect 17007 14660 17013 14662
rect 16705 14651 17013 14660
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16040 12850 16068 13262
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15580 11694 15608 12786
rect 16040 12238 16068 12786
rect 16408 12714 16436 13262
rect 16500 12782 16528 13670
rect 16592 13308 16620 14486
rect 17052 13954 17080 14878
rect 17236 14618 17264 15438
rect 17696 15366 17724 16102
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 15706 17816 15982
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 18064 15502 18092 16458
rect 18156 15586 18184 17750
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18248 17338 18276 17546
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17338 18460 17478
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18524 16726 18552 16934
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 19076 16182 19104 20402
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19168 19446 19196 19790
rect 19352 19530 19380 26930
rect 23007 26684 23315 26693
rect 23007 26682 23013 26684
rect 23069 26682 23093 26684
rect 23149 26682 23173 26684
rect 23229 26682 23253 26684
rect 23309 26682 23315 26684
rect 23069 26630 23071 26682
rect 23251 26630 23253 26682
rect 23007 26628 23013 26630
rect 23069 26628 23093 26630
rect 23149 26628 23173 26630
rect 23229 26628 23253 26630
rect 23309 26628 23315 26630
rect 23007 26619 23315 26628
rect 20720 26444 20772 26450
rect 20720 26386 20772 26392
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19444 25362 19472 25842
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19444 22506 19472 25298
rect 19708 25220 19760 25226
rect 19708 25162 19760 25168
rect 19720 24954 19748 25162
rect 20088 24954 20116 25774
rect 20732 25226 20760 26386
rect 20812 26308 20864 26314
rect 20812 26250 20864 26256
rect 20824 25974 20852 26250
rect 23400 26042 23428 26930
rect 23667 26140 23975 26149
rect 23667 26138 23673 26140
rect 23729 26138 23753 26140
rect 23809 26138 23833 26140
rect 23889 26138 23913 26140
rect 23969 26138 23975 26140
rect 23729 26086 23731 26138
rect 23911 26086 23913 26138
rect 23667 26084 23673 26086
rect 23729 26084 23753 26086
rect 23809 26084 23833 26086
rect 23889 26084 23913 26086
rect 23969 26084 23975 26086
rect 23667 26075 23975 26084
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 20812 25968 20864 25974
rect 20812 25910 20864 25916
rect 23572 25968 23624 25974
rect 23572 25910 23624 25916
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 20812 25424 20864 25430
rect 20812 25366 20864 25372
rect 20720 25220 20772 25226
rect 20720 25162 20772 25168
rect 20824 24970 20852 25366
rect 21284 25294 21312 25638
rect 21364 25356 21416 25362
rect 21416 25316 21496 25344
rect 21364 25298 21416 25304
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 19708 24948 19760 24954
rect 19708 24890 19760 24896
rect 20076 24948 20128 24954
rect 20076 24890 20128 24896
rect 20732 24942 20852 24970
rect 20732 24886 20760 24942
rect 20720 24880 20772 24886
rect 20720 24822 20772 24828
rect 21192 24818 21220 25094
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 20076 24744 20128 24750
rect 20076 24686 20128 24692
rect 19904 24070 19932 24686
rect 20088 24206 20116 24686
rect 20548 24342 20576 24754
rect 20640 24392 20668 24754
rect 20824 24614 20852 24754
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 20720 24404 20772 24410
rect 20640 24364 20720 24392
rect 20720 24346 20772 24352
rect 20536 24336 20588 24342
rect 20536 24278 20588 24284
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20258 24168 20314 24177
rect 20824 24138 20852 24550
rect 21192 24410 21220 24754
rect 21284 24682 21312 25230
rect 21364 25220 21416 25226
rect 21364 25162 21416 25168
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20258 24103 20314 24112
rect 20720 24132 20772 24138
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19628 22658 19656 23258
rect 19800 23248 19852 23254
rect 19800 23190 19852 23196
rect 20074 23216 20130 23225
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19720 22778 19748 23054
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19812 22710 19840 23190
rect 20074 23151 20076 23160
rect 20128 23151 20130 23160
rect 20076 23122 20128 23128
rect 20272 23120 20300 24103
rect 20720 24074 20772 24080
rect 20812 24132 20864 24138
rect 20812 24074 20864 24080
rect 20732 23526 20760 24074
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20350 23352 20406 23361
rect 20350 23287 20406 23296
rect 20168 23112 20220 23118
rect 19890 23080 19946 23089
rect 19890 23015 19892 23024
rect 19944 23015 19946 23024
rect 20088 23060 20168 23066
rect 20088 23054 20220 23060
rect 20260 23114 20312 23120
rect 20260 23056 20312 23062
rect 20088 23038 20208 23054
rect 19892 22986 19944 22992
rect 20088 22778 20116 23038
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 19800 22704 19852 22710
rect 19536 22642 19748 22658
rect 19800 22646 19852 22652
rect 19536 22636 19760 22642
rect 19536 22630 19708 22636
rect 19432 22500 19484 22506
rect 19432 22442 19484 22448
rect 19536 22030 19564 22630
rect 19708 22578 19760 22584
rect 19616 22568 19668 22574
rect 19616 22510 19668 22516
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19628 21010 19656 22510
rect 19708 22432 19760 22438
rect 19708 22374 19760 22380
rect 19720 21962 19748 22374
rect 19812 22098 19840 22646
rect 20088 22234 20116 22714
rect 20364 22574 20392 23287
rect 20456 23118 20484 23462
rect 20718 23352 20774 23361
rect 20628 23316 20680 23322
rect 20718 23287 20720 23296
rect 20628 23258 20680 23264
rect 20772 23287 20774 23296
rect 20720 23258 20772 23264
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20640 22964 20668 23258
rect 20718 23216 20774 23225
rect 20718 23151 20720 23160
rect 20772 23151 20774 23160
rect 20720 23122 20772 23128
rect 20824 23118 20852 24074
rect 20916 23866 20944 24210
rect 21088 24200 21140 24206
rect 21192 24188 21220 24346
rect 21140 24160 21220 24188
rect 21088 24142 21140 24148
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 21192 23798 21220 24160
rect 21180 23792 21232 23798
rect 21180 23734 21232 23740
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 21008 23322 21036 23666
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20904 22976 20956 22982
rect 20640 22936 20904 22964
rect 20904 22918 20956 22924
rect 21008 22574 21036 23122
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 21100 22438 21128 23054
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19800 22092 19852 22098
rect 21192 22094 21220 23734
rect 21284 23526 21312 24618
rect 21376 24206 21404 25162
rect 21468 24682 21496 25316
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 21824 25152 21876 25158
rect 21824 25094 21876 25100
rect 21836 24886 21864 25094
rect 21824 24880 21876 24886
rect 21824 24822 21876 24828
rect 22020 24834 22048 25230
rect 22112 25158 22140 25842
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22480 24954 22508 25230
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 22020 24818 22140 24834
rect 22204 24818 22232 24890
rect 22480 24818 22508 24890
rect 22020 24812 22152 24818
rect 22020 24806 22100 24812
rect 22100 24754 22152 24760
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 21456 24676 21508 24682
rect 21456 24618 21508 24624
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21376 24070 21404 24142
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21376 23798 21404 24006
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21376 23254 21404 23734
rect 21364 23248 21416 23254
rect 21364 23190 21416 23196
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21284 23089 21312 23122
rect 21270 23080 21326 23089
rect 21270 23015 21326 23024
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21376 22506 21404 22918
rect 21468 22778 21496 24618
rect 22388 24410 22416 24754
rect 22572 24410 22600 25774
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22204 23730 22232 24210
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22296 23798 22324 24142
rect 22572 23866 22600 24346
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22284 23792 22336 23798
rect 22284 23734 22336 23740
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22572 23322 22600 23666
rect 22664 23662 22692 25842
rect 23007 25596 23315 25605
rect 23007 25594 23013 25596
rect 23069 25594 23093 25596
rect 23149 25594 23173 25596
rect 23229 25594 23253 25596
rect 23309 25594 23315 25596
rect 23069 25542 23071 25594
rect 23251 25542 23253 25594
rect 23007 25540 23013 25542
rect 23069 25540 23093 25542
rect 23149 25540 23173 25542
rect 23229 25540 23253 25542
rect 23309 25540 23315 25542
rect 23007 25531 23315 25540
rect 23584 25498 23612 25910
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 24412 25294 24440 25638
rect 24308 25288 24360 25294
rect 24308 25230 24360 25236
rect 24400 25288 24452 25294
rect 25780 25288 25832 25294
rect 24400 25230 24452 25236
rect 25778 25256 25780 25265
rect 25832 25256 25834 25265
rect 22744 25152 22796 25158
rect 22744 25094 22796 25100
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22376 23248 22428 23254
rect 22296 23208 22376 23236
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21548 22704 21600 22710
rect 21548 22646 21600 22652
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21560 22098 21588 22646
rect 22296 22574 22324 23208
rect 22376 23190 22428 23196
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22572 22778 22600 22986
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22664 22642 22692 23598
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 19800 22034 19852 22040
rect 21100 22066 21220 22094
rect 21548 22092 21600 22098
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19720 21146 19748 21898
rect 19812 21350 19840 22034
rect 21100 21894 21128 22066
rect 21548 22034 21600 22040
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19430 20904 19486 20913
rect 19430 20839 19486 20848
rect 19444 19922 19472 20839
rect 19628 20602 19656 20946
rect 19892 20868 19944 20874
rect 19892 20810 19944 20816
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 19904 20058 19932 20810
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19260 19502 19380 19530
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 18248 15706 18276 16118
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 19076 15638 19104 16118
rect 19064 15632 19116 15638
rect 18156 15558 18276 15586
rect 19064 15574 19116 15580
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17365 15260 17673 15269
rect 17365 15258 17371 15260
rect 17427 15258 17451 15260
rect 17507 15258 17531 15260
rect 17587 15258 17611 15260
rect 17667 15258 17673 15260
rect 17427 15206 17429 15258
rect 17609 15206 17611 15258
rect 17365 15204 17371 15206
rect 17427 15204 17451 15206
rect 17507 15204 17531 15206
rect 17587 15204 17611 15206
rect 17667 15204 17673 15206
rect 17365 15195 17673 15204
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17328 14414 17356 14962
rect 17880 14550 17908 15370
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17144 14074 17172 14350
rect 17365 14172 17673 14181
rect 17365 14170 17371 14172
rect 17427 14170 17451 14172
rect 17507 14170 17531 14172
rect 17587 14170 17611 14172
rect 17667 14170 17673 14172
rect 17427 14118 17429 14170
rect 17609 14118 17611 14170
rect 17365 14116 17371 14118
rect 17427 14116 17451 14118
rect 17507 14116 17531 14118
rect 17587 14116 17611 14118
rect 17667 14116 17673 14118
rect 17365 14107 17673 14116
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17224 14000 17276 14006
rect 16960 13948 17224 13954
rect 16960 13942 17276 13948
rect 16960 13926 17264 13942
rect 16960 13870 16988 13926
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 16705 13628 17013 13637
rect 16705 13626 16711 13628
rect 16767 13626 16791 13628
rect 16847 13626 16871 13628
rect 16927 13626 16951 13628
rect 17007 13626 17013 13628
rect 16767 13574 16769 13626
rect 16949 13574 16951 13626
rect 16705 13572 16711 13574
rect 16767 13572 16791 13574
rect 16847 13572 16871 13574
rect 16927 13572 16951 13574
rect 17007 13572 17013 13574
rect 16705 13563 17013 13572
rect 16672 13320 16724 13326
rect 16592 13280 16672 13308
rect 16672 13262 16724 13268
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16408 12374 16436 12650
rect 16500 12424 16528 12718
rect 16705 12540 17013 12549
rect 16705 12538 16711 12540
rect 16767 12538 16791 12540
rect 16847 12538 16871 12540
rect 16927 12538 16951 12540
rect 17007 12538 17013 12540
rect 16767 12486 16769 12538
rect 16949 12486 16951 12538
rect 16705 12484 16711 12486
rect 16767 12484 16791 12486
rect 16847 12484 16871 12486
rect 16927 12484 16951 12486
rect 17007 12484 17013 12486
rect 16705 12475 17013 12484
rect 17052 12442 17080 13262
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 16672 12436 16724 12442
rect 16500 12396 16672 12424
rect 16672 12378 16724 12384
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15580 11150 15608 11630
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15672 11354 15700 11562
rect 16040 11558 16068 12174
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15580 10674 15608 11086
rect 16040 11082 16068 11494
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 15304 9382 15332 10542
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15106 9072 15162 9081
rect 14832 9036 14884 9042
rect 15106 9007 15162 9016
rect 14832 8978 14884 8984
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14752 5914 14780 6326
rect 15028 6322 15056 6598
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15120 6118 15148 6938
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14752 5030 14780 5510
rect 14936 5234 14964 5510
rect 15120 5302 15148 6054
rect 15212 5370 15240 8910
rect 15304 8498 15332 9318
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 15304 6798 15332 7414
rect 15396 7002 15424 9590
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15488 7834 15516 8026
rect 15488 7806 15608 7834
rect 15672 7818 15700 10134
rect 15764 8906 15792 10406
rect 16316 9994 16344 10542
rect 16408 10062 16436 12310
rect 17144 11830 17172 13126
rect 17236 12782 17264 13806
rect 17512 13326 17540 14010
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17604 13190 17632 13942
rect 17880 13920 17908 14486
rect 17788 13892 17908 13920
rect 17788 13530 17816 13892
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17880 13394 17908 13738
rect 17972 13530 18000 14758
rect 18064 14006 18092 14962
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18156 14618 18184 14894
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18156 14414 18184 14554
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17365 13084 17673 13093
rect 17365 13082 17371 13084
rect 17427 13082 17451 13084
rect 17507 13082 17531 13084
rect 17587 13082 17611 13084
rect 17667 13082 17673 13084
rect 17427 13030 17429 13082
rect 17609 13030 17611 13082
rect 17365 13028 17371 13030
rect 17427 13028 17451 13030
rect 17507 13028 17531 13030
rect 17587 13028 17611 13030
rect 17667 13028 17673 13030
rect 17365 13019 17673 13028
rect 17788 12986 17816 13262
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17328 12374 17356 12786
rect 17776 12640 17828 12646
rect 17880 12628 17908 13330
rect 17972 13258 18000 13466
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17828 12600 17908 12628
rect 17776 12582 17828 12588
rect 17316 12368 17368 12374
rect 17236 12328 17316 12356
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 16705 11452 17013 11461
rect 16705 11450 16711 11452
rect 16767 11450 16791 11452
rect 16847 11450 16871 11452
rect 16927 11450 16951 11452
rect 17007 11450 17013 11452
rect 16767 11398 16769 11450
rect 16949 11398 16951 11450
rect 16705 11396 16711 11398
rect 16767 11396 16791 11398
rect 16847 11396 16871 11398
rect 16927 11396 16951 11398
rect 17007 11396 17013 11398
rect 16705 11387 17013 11396
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9654 16160 9862
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16316 9602 16344 9930
rect 16212 9580 16264 9586
rect 16316 9574 16436 9602
rect 16212 9522 16264 9528
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 16224 8498 16252 9522
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16316 8634 16344 9454
rect 16408 9450 16436 9574
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16396 9172 16448 9178
rect 16592 9160 16620 11222
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16705 10364 17013 10373
rect 16705 10362 16711 10364
rect 16767 10362 16791 10364
rect 16847 10362 16871 10364
rect 16927 10362 16951 10364
rect 17007 10362 17013 10364
rect 16767 10310 16769 10362
rect 16949 10310 16951 10362
rect 16705 10308 16711 10310
rect 16767 10308 16791 10310
rect 16847 10308 16871 10310
rect 16927 10308 16951 10310
rect 17007 10308 17013 10310
rect 16705 10299 17013 10308
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16684 9654 16712 9998
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16960 9450 16988 10202
rect 17052 10198 17080 11018
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16705 9276 17013 9285
rect 16705 9274 16711 9276
rect 16767 9274 16791 9276
rect 16847 9274 16871 9276
rect 16927 9274 16951 9276
rect 17007 9274 17013 9276
rect 16767 9222 16769 9274
rect 16949 9222 16951 9274
rect 16705 9220 16711 9222
rect 16767 9220 16791 9222
rect 16847 9220 16871 9222
rect 16927 9220 16951 9222
rect 17007 9220 17013 9222
rect 16705 9211 17013 9220
rect 17144 9178 17172 9862
rect 17236 9654 17264 12328
rect 17316 12310 17368 12316
rect 17788 12238 17816 12582
rect 17972 12458 18000 12922
rect 18064 12918 18092 13126
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17880 12430 18000 12458
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17365 11996 17673 12005
rect 17365 11994 17371 11996
rect 17427 11994 17451 11996
rect 17507 11994 17531 11996
rect 17587 11994 17611 11996
rect 17667 11994 17673 11996
rect 17427 11942 17429 11994
rect 17609 11942 17611 11994
rect 17365 11940 17371 11942
rect 17427 11940 17451 11942
rect 17507 11940 17531 11942
rect 17587 11940 17611 11942
rect 17667 11940 17673 11942
rect 17365 11931 17673 11940
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17788 11354 17816 11766
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17365 10908 17673 10917
rect 17365 10906 17371 10908
rect 17427 10906 17451 10908
rect 17507 10906 17531 10908
rect 17587 10906 17611 10908
rect 17667 10906 17673 10908
rect 17427 10854 17429 10906
rect 17609 10854 17611 10906
rect 17365 10852 17371 10854
rect 17427 10852 17451 10854
rect 17507 10852 17531 10854
rect 17587 10852 17611 10854
rect 17667 10852 17673 10854
rect 17365 10843 17673 10852
rect 17365 9820 17673 9829
rect 17365 9818 17371 9820
rect 17427 9818 17451 9820
rect 17507 9818 17531 9820
rect 17587 9818 17611 9820
rect 17667 9818 17673 9820
rect 17427 9766 17429 9818
rect 17609 9766 17611 9818
rect 17365 9764 17371 9766
rect 17427 9764 17451 9766
rect 17507 9764 17531 9766
rect 17587 9764 17611 9766
rect 17667 9764 17673 9766
rect 17365 9755 17673 9764
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17880 9568 17908 12430
rect 18064 11218 18092 12854
rect 18156 12714 18184 14350
rect 18248 12986 18276 15558
rect 19168 15502 19196 19382
rect 19260 18970 19288 19502
rect 19996 19446 20024 21422
rect 21376 21146 21404 21422
rect 21364 21140 21416 21146
rect 21284 21100 21364 21128
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 19922 20484 20402
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20180 19446 20208 19790
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19352 18970 19380 19314
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20088 18834 20116 18906
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19628 17678 19656 18702
rect 19812 18630 19840 18702
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19720 17542 19748 18362
rect 19812 18358 19840 18566
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19812 17202 19840 18022
rect 20088 17746 20116 18770
rect 20180 18426 20208 19382
rect 20456 19242 20484 19722
rect 20548 19514 20576 19790
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20640 19258 20668 20334
rect 20916 19802 20944 20334
rect 21284 20262 21312 21100
rect 21364 21082 21416 21088
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 20996 20256 21048 20262
rect 21272 20256 21324 20262
rect 20996 20198 21048 20204
rect 21100 20216 21272 20244
rect 21008 19922 21036 20198
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20916 19774 21036 19802
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20916 19446 20944 19654
rect 20720 19440 20772 19446
rect 20904 19440 20956 19446
rect 20772 19400 20852 19428
rect 20720 19382 20772 19388
rect 20720 19304 20772 19310
rect 20640 19252 20720 19258
rect 20640 19246 20772 19252
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20640 19230 20760 19246
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20272 18086 20300 18906
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18358 20392 18566
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20456 18154 20484 19178
rect 20640 18970 20668 19230
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20444 18148 20496 18154
rect 20444 18090 20496 18096
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19904 16658 19932 17614
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19996 17134 20024 17546
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 20088 17066 20116 17478
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 20088 16946 20116 17002
rect 20088 16918 20208 16946
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 20180 16522 20208 16918
rect 20272 16697 20300 17682
rect 20548 17678 20576 18634
rect 20640 18222 20668 18906
rect 20732 18766 20760 18906
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20824 18306 20852 19400
rect 20904 19382 20956 19388
rect 20732 18290 20852 18306
rect 21008 18290 21036 19774
rect 21100 19378 21128 20216
rect 21272 20198 21324 20204
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 19854 21404 20198
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21100 18834 21128 18906
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 21100 18290 21128 18566
rect 20720 18284 20852 18290
rect 20772 18278 20852 18284
rect 20996 18284 21048 18290
rect 20720 18226 20772 18232
rect 20996 18226 21048 18232
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20732 17610 20760 18226
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20258 16688 20314 16697
rect 20258 16623 20314 16632
rect 20272 16590 20300 16623
rect 20548 16590 20576 17070
rect 20732 16794 20760 17546
rect 21008 17134 21036 18090
rect 21192 17678 21220 19722
rect 21284 19514 21312 19790
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21468 19242 21496 20402
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21560 19174 21588 19722
rect 21652 19446 21680 20334
rect 21824 19984 21876 19990
rect 21824 19926 21876 19932
rect 21640 19440 21692 19446
rect 21640 19382 21692 19388
rect 21836 19378 21864 19926
rect 22020 19922 22048 20470
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22296 19394 22324 19858
rect 22020 19378 22324 19394
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 22008 19372 22324 19378
rect 22060 19366 22324 19372
rect 22008 19314 22060 19320
rect 22020 19242 22048 19314
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16794 20944 16934
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20812 16720 20864 16726
rect 21008 16674 21036 17070
rect 20812 16662 20864 16668
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20536 16584 20588 16590
rect 20720 16584 20772 16590
rect 20536 16526 20588 16532
rect 20718 16552 20720 16561
rect 20772 16552 20774 16561
rect 20168 16516 20220 16522
rect 20718 16487 20774 16496
rect 20168 16458 20220 16464
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18340 13326 18368 14826
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14414 18552 14758
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18708 14090 18736 14350
rect 18708 14062 18828 14090
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18708 13326 18736 13942
rect 18800 13326 18828 14062
rect 18892 13802 18920 14962
rect 19260 14482 19288 16186
rect 20732 15586 20760 16186
rect 20824 16114 20852 16662
rect 20916 16646 21036 16674
rect 20916 16402 20944 16646
rect 21192 16538 21220 17614
rect 21284 17338 21312 18702
rect 21376 18426 21404 18702
rect 21560 18698 21588 19110
rect 22756 18873 22784 25094
rect 23007 24508 23315 24517
rect 23007 24506 23013 24508
rect 23069 24506 23093 24508
rect 23149 24506 23173 24508
rect 23229 24506 23253 24508
rect 23309 24506 23315 24508
rect 23069 24454 23071 24506
rect 23251 24454 23253 24506
rect 23007 24452 23013 24454
rect 23069 24452 23093 24454
rect 23149 24452 23173 24454
rect 23229 24452 23253 24454
rect 23309 24452 23315 24454
rect 23007 24443 23315 24452
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23112 24200 23164 24206
rect 23110 24168 23112 24177
rect 23164 24168 23166 24177
rect 22928 24132 22980 24138
rect 23110 24103 23166 24112
rect 22928 24074 22980 24080
rect 22940 23866 22968 24074
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 23400 23526 23428 24346
rect 23492 24342 23520 25094
rect 23667 25052 23975 25061
rect 23667 25050 23673 25052
rect 23729 25050 23753 25052
rect 23809 25050 23833 25052
rect 23889 25050 23913 25052
rect 23969 25050 23975 25052
rect 23729 24998 23731 25050
rect 23911 24998 23913 25050
rect 23667 24996 23673 24998
rect 23729 24996 23753 24998
rect 23809 24996 23833 24998
rect 23889 24996 23913 24998
rect 23969 24996 23975 24998
rect 23667 24987 23975 24996
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 24320 24206 24348 25230
rect 25778 25191 25834 25200
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 25228 25152 25280 25158
rect 25228 25094 25280 25100
rect 23572 24200 23624 24206
rect 24308 24200 24360 24206
rect 23572 24142 23624 24148
rect 23754 24168 23810 24177
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23730 23520 24006
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 22940 22642 22968 23462
rect 23007 23420 23315 23429
rect 23007 23418 23013 23420
rect 23069 23418 23093 23420
rect 23149 23418 23173 23420
rect 23229 23418 23253 23420
rect 23309 23418 23315 23420
rect 23069 23366 23071 23418
rect 23251 23366 23253 23418
rect 23007 23364 23013 23366
rect 23069 23364 23093 23366
rect 23149 23364 23173 23366
rect 23229 23364 23253 23366
rect 23309 23364 23315 23366
rect 23007 23355 23315 23364
rect 23400 23322 23428 23462
rect 23584 23322 23612 24142
rect 24308 24142 24360 24148
rect 23754 24103 23756 24112
rect 23808 24103 23810 24112
rect 23756 24074 23808 24080
rect 23667 23964 23975 23973
rect 23667 23962 23673 23964
rect 23729 23962 23753 23964
rect 23809 23962 23833 23964
rect 23889 23962 23913 23964
rect 23969 23962 23975 23964
rect 23729 23910 23731 23962
rect 23911 23910 23913 23962
rect 23667 23908 23673 23910
rect 23729 23908 23753 23910
rect 23809 23908 23833 23910
rect 23889 23908 23913 23910
rect 23969 23908 23975 23910
rect 23667 23899 23975 23908
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23676 23118 23704 23462
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23848 23112 23900 23118
rect 24216 23112 24268 23118
rect 23900 23072 24072 23100
rect 23848 23054 23900 23060
rect 23667 22876 23975 22885
rect 23667 22874 23673 22876
rect 23729 22874 23753 22876
rect 23809 22874 23833 22876
rect 23889 22874 23913 22876
rect 23969 22874 23975 22876
rect 23729 22822 23731 22874
rect 23911 22822 23913 22874
rect 23667 22820 23673 22822
rect 23729 22820 23753 22822
rect 23809 22820 23833 22822
rect 23889 22820 23913 22822
rect 23969 22820 23975 22822
rect 23667 22811 23975 22820
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 23007 22332 23315 22341
rect 23007 22330 23013 22332
rect 23069 22330 23093 22332
rect 23149 22330 23173 22332
rect 23229 22330 23253 22332
rect 23309 22330 23315 22332
rect 23069 22278 23071 22330
rect 23251 22278 23253 22330
rect 23007 22276 23013 22278
rect 23069 22276 23093 22278
rect 23149 22276 23173 22278
rect 23229 22276 23253 22278
rect 23309 22276 23315 22278
rect 23007 22267 23315 22276
rect 23768 22098 23796 22646
rect 24044 22574 24072 23072
rect 24216 23054 24268 23060
rect 24228 22710 24256 23054
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23667 21788 23975 21797
rect 23667 21786 23673 21788
rect 23729 21786 23753 21788
rect 23809 21786 23833 21788
rect 23889 21786 23913 21788
rect 23969 21786 23975 21788
rect 23729 21734 23731 21786
rect 23911 21734 23913 21786
rect 23667 21732 23673 21734
rect 23729 21732 23753 21734
rect 23809 21732 23833 21734
rect 23889 21732 23913 21734
rect 23969 21732 23975 21734
rect 23667 21723 23975 21732
rect 23007 21244 23315 21253
rect 23007 21242 23013 21244
rect 23069 21242 23093 21244
rect 23149 21242 23173 21244
rect 23229 21242 23253 21244
rect 23309 21242 23315 21244
rect 23069 21190 23071 21242
rect 23251 21190 23253 21242
rect 23007 21188 23013 21190
rect 23069 21188 23093 21190
rect 23149 21188 23173 21190
rect 23229 21188 23253 21190
rect 23309 21188 23315 21190
rect 23007 21179 23315 21188
rect 24044 21010 24072 22510
rect 24320 22030 24348 24142
rect 25056 24138 25084 25094
rect 25044 24132 25096 24138
rect 25044 24074 25096 24080
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24504 23798 24532 24006
rect 24492 23792 24544 23798
rect 24492 23734 24544 23740
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24320 20942 24348 21966
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 23400 20466 23428 20742
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23007 20156 23315 20165
rect 23007 20154 23013 20156
rect 23069 20154 23093 20156
rect 23149 20154 23173 20156
rect 23229 20154 23253 20156
rect 23309 20154 23315 20156
rect 23069 20102 23071 20154
rect 23251 20102 23253 20154
rect 23007 20100 23013 20102
rect 23069 20100 23093 20102
rect 23149 20100 23173 20102
rect 23229 20100 23253 20102
rect 23309 20100 23315 20102
rect 23007 20091 23315 20100
rect 23296 19780 23348 19786
rect 23296 19722 23348 19728
rect 23308 19514 23336 19722
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23492 19394 23520 20878
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 23667 20700 23975 20709
rect 23667 20698 23673 20700
rect 23729 20698 23753 20700
rect 23809 20698 23833 20700
rect 23889 20698 23913 20700
rect 23969 20698 23975 20700
rect 23729 20646 23731 20698
rect 23911 20646 23913 20698
rect 23667 20644 23673 20646
rect 23729 20644 23753 20646
rect 23809 20644 23833 20646
rect 23889 20644 23913 20646
rect 23969 20644 23975 20646
rect 23667 20635 23975 20644
rect 24044 20534 24072 20742
rect 24780 20534 24808 20878
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 24768 20528 24820 20534
rect 24768 20470 24820 20476
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 23667 19612 23975 19621
rect 23667 19610 23673 19612
rect 23729 19610 23753 19612
rect 23809 19610 23833 19612
rect 23889 19610 23913 19612
rect 23969 19610 23975 19612
rect 23729 19558 23731 19610
rect 23911 19558 23913 19610
rect 23667 19556 23673 19558
rect 23729 19556 23753 19558
rect 23809 19556 23833 19558
rect 23889 19556 23913 19558
rect 23969 19556 23975 19558
rect 23667 19547 23975 19556
rect 23400 19378 23520 19394
rect 23388 19372 23520 19378
rect 23440 19366 23520 19372
rect 23388 19314 23440 19320
rect 23007 19068 23315 19077
rect 23007 19066 23013 19068
rect 23069 19066 23093 19068
rect 23149 19066 23173 19068
rect 23229 19066 23253 19068
rect 23309 19066 23315 19068
rect 23069 19014 23071 19066
rect 23251 19014 23253 19066
rect 23007 19012 23013 19014
rect 23069 19012 23093 19014
rect 23149 19012 23173 19014
rect 23229 19012 23253 19014
rect 23309 19012 23315 19014
rect 23007 19003 23315 19012
rect 23492 18902 23520 19366
rect 23480 18896 23532 18902
rect 22742 18864 22798 18873
rect 23480 18838 23532 18844
rect 22742 18799 22798 18808
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 21456 18692 21508 18698
rect 21456 18634 21508 18640
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21468 18358 21496 18634
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21560 17898 21588 18634
rect 21376 17870 21588 17898
rect 21376 17610 21404 17870
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21376 16658 21404 17546
rect 21468 17202 21496 17614
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 22008 17196 22060 17202
rect 22112 17184 22140 18702
rect 23007 17980 23315 17989
rect 23007 17978 23013 17980
rect 23069 17978 23093 17980
rect 23149 17978 23173 17980
rect 23229 17978 23253 17980
rect 23309 17978 23315 17980
rect 23069 17926 23071 17978
rect 23251 17926 23253 17978
rect 23007 17924 23013 17926
rect 23069 17924 23093 17926
rect 23149 17924 23173 17926
rect 23229 17924 23253 17926
rect 23309 17924 23315 17926
rect 23007 17915 23315 17924
rect 23492 17746 23520 18838
rect 23667 18524 23975 18533
rect 23667 18522 23673 18524
rect 23729 18522 23753 18524
rect 23809 18522 23833 18524
rect 23889 18522 23913 18524
rect 23969 18522 23975 18524
rect 23729 18470 23731 18522
rect 23911 18470 23913 18522
rect 23667 18468 23673 18470
rect 23729 18468 23753 18470
rect 23809 18468 23833 18470
rect 23889 18468 23913 18470
rect 23969 18468 23975 18470
rect 23667 18459 23975 18468
rect 25148 18426 25176 20334
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25240 18329 25268 25094
rect 27080 23769 27108 28825
rect 27066 23760 27122 23769
rect 27066 23695 27122 23704
rect 25780 21548 25832 21554
rect 25780 21490 25832 21496
rect 25792 21185 25820 21490
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25778 21176 25834 21185
rect 25778 21111 25834 21120
rect 25976 20058 26004 21286
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 25226 18320 25282 18329
rect 25044 18284 25096 18290
rect 25226 18255 25282 18264
rect 25044 18226 25096 18232
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22296 17270 22324 17478
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22060 17156 22140 17184
rect 22008 17138 22060 17144
rect 22112 16658 22140 17156
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 21272 16584 21324 16590
rect 21008 16522 21220 16538
rect 20996 16516 21220 16522
rect 21048 16510 21220 16516
rect 20996 16458 21048 16464
rect 21088 16448 21140 16454
rect 20916 16374 21036 16402
rect 21088 16390 21140 16396
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20640 15570 20760 15586
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 20628 15564 20760 15570
rect 20680 15558 20760 15564
rect 20628 15506 20680 15512
rect 19996 15026 20024 15506
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 19248 14476 19300 14482
rect 19168 14436 19248 14464
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18984 14074 19012 14350
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 19168 13938 19196 14436
rect 19248 14418 19300 14424
rect 20088 14346 20116 14758
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18892 13462 18920 13738
rect 19444 13462 19472 14282
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19812 13530 19840 13806
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 18892 13326 18920 13398
rect 20180 13326 20208 14214
rect 20272 14006 20300 14758
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 13530 20392 13670
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18880 13320 18932 13326
rect 19064 13320 19116 13326
rect 18932 13280 19064 13308
rect 18880 13262 18932 13268
rect 19064 13262 19116 13268
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18616 12986 18644 13126
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18892 12850 18920 13262
rect 20364 12850 20392 13466
rect 20732 13394 20760 15558
rect 20824 15502 20852 16050
rect 21008 16046 21036 16374
rect 21100 16182 21128 16390
rect 21192 16250 21220 16510
rect 21270 16552 21272 16561
rect 21324 16552 21326 16561
rect 21270 16487 21326 16496
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 21284 16046 21312 16487
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21008 15706 21036 15982
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21468 15570 21496 16594
rect 22756 16522 22784 17478
rect 23007 16892 23315 16901
rect 23007 16890 23013 16892
rect 23069 16890 23093 16892
rect 23149 16890 23173 16892
rect 23229 16890 23253 16892
rect 23309 16890 23315 16892
rect 23069 16838 23071 16890
rect 23251 16838 23253 16890
rect 23007 16836 23013 16838
rect 23069 16836 23093 16838
rect 23149 16836 23173 16838
rect 23229 16836 23253 16838
rect 23309 16836 23315 16838
rect 23007 16827 23315 16836
rect 23204 16720 23256 16726
rect 23202 16688 23204 16697
rect 23256 16688 23258 16697
rect 23202 16623 23258 16632
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 21836 15978 21864 16458
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 23007 15804 23315 15813
rect 23007 15802 23013 15804
rect 23069 15802 23093 15804
rect 23149 15802 23173 15804
rect 23229 15802 23253 15804
rect 23309 15802 23315 15804
rect 23069 15750 23071 15802
rect 23251 15750 23253 15802
rect 23007 15748 23013 15750
rect 23069 15748 23093 15750
rect 23149 15748 23173 15750
rect 23229 15748 23253 15750
rect 23309 15748 23315 15750
rect 23007 15739 23315 15748
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21100 15162 21128 15370
rect 23400 15366 23428 17614
rect 23492 17218 23520 17682
rect 23667 17436 23975 17445
rect 23667 17434 23673 17436
rect 23729 17434 23753 17436
rect 23809 17434 23833 17436
rect 23889 17434 23913 17436
rect 23969 17434 23975 17436
rect 23729 17382 23731 17434
rect 23911 17382 23913 17434
rect 23667 17380 23673 17382
rect 23729 17380 23753 17382
rect 23809 17380 23833 17382
rect 23889 17380 23913 17382
rect 23969 17380 23975 17382
rect 23667 17371 23975 17380
rect 23492 17190 23612 17218
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23492 16454 23520 17070
rect 23584 16658 23612 17190
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23667 16348 23975 16357
rect 23667 16346 23673 16348
rect 23729 16346 23753 16348
rect 23809 16346 23833 16348
rect 23889 16346 23913 16348
rect 23969 16346 23975 16348
rect 23729 16294 23731 16346
rect 23911 16294 23913 16346
rect 23667 16292 23673 16294
rect 23729 16292 23753 16294
rect 23809 16292 23833 16294
rect 23889 16292 23913 16294
rect 23969 16292 23975 16294
rect 23667 16283 23975 16292
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 23667 15260 23975 15269
rect 23667 15258 23673 15260
rect 23729 15258 23753 15260
rect 23809 15258 23833 15260
rect 23889 15258 23913 15260
rect 23969 15258 23975 15260
rect 23729 15206 23731 15258
rect 23911 15206 23913 15258
rect 23667 15204 23673 15206
rect 23729 15204 23753 15206
rect 23809 15204 23833 15206
rect 23889 15204 23913 15206
rect 23969 15204 23975 15206
rect 23667 15195 23975 15204
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 23007 14716 23315 14725
rect 23007 14714 23013 14716
rect 23069 14714 23093 14716
rect 23149 14714 23173 14716
rect 23229 14714 23253 14716
rect 23309 14714 23315 14716
rect 23069 14662 23071 14714
rect 23251 14662 23253 14714
rect 23007 14660 23013 14662
rect 23069 14660 23093 14662
rect 23149 14660 23173 14662
rect 23229 14660 23253 14662
rect 23309 14660 23315 14662
rect 23007 14651 23315 14660
rect 23667 14172 23975 14181
rect 23667 14170 23673 14172
rect 23729 14170 23753 14172
rect 23809 14170 23833 14172
rect 23889 14170 23913 14172
rect 23969 14170 23975 14172
rect 23729 14118 23731 14170
rect 23911 14118 23913 14170
rect 23667 14116 23673 14118
rect 23729 14116 23753 14118
rect 23809 14116 23833 14118
rect 23889 14116 23913 14118
rect 23969 14116 23975 14118
rect 23667 14107 23975 14116
rect 23007 13628 23315 13637
rect 23007 13626 23013 13628
rect 23069 13626 23093 13628
rect 23149 13626 23173 13628
rect 23229 13626 23253 13628
rect 23309 13626 23315 13628
rect 23069 13574 23071 13626
rect 23251 13574 23253 13626
rect 23007 13572 23013 13574
rect 23069 13572 23093 13574
rect 23149 13572 23173 13574
rect 23229 13572 23253 13574
rect 23309 13572 23315 13574
rect 23007 13563 23315 13572
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 21100 12986 21128 13194
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18248 12170 18276 12718
rect 18892 12434 18920 12786
rect 21192 12434 21220 12786
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 18800 12406 18920 12434
rect 21008 12406 21220 12434
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18248 11558 18276 12106
rect 18800 11898 18828 12406
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18420 11824 18472 11830
rect 20732 11801 20760 12174
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20916 11898 20944 12106
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 18420 11766 18472 11772
rect 20718 11792 20774 11801
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17972 10810 18000 11154
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17788 9540 17908 9568
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17512 9178 17540 9318
rect 17132 9172 17184 9178
rect 16592 9132 16712 9160
rect 16396 9114 16448 9120
rect 16408 8634 16436 9114
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16500 8566 16528 8774
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 15580 7750 15608 7806
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6254 15332 6734
rect 15488 6662 15516 7686
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 6322 15516 6598
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15304 5794 15332 6190
rect 15580 5914 15608 6666
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15304 5766 15424 5794
rect 15396 5710 15424 5766
rect 15672 5710 15700 7754
rect 16132 7290 16160 8230
rect 16224 8090 16252 8230
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16500 8022 16528 8502
rect 16592 8090 16620 8978
rect 16684 8566 16712 9132
rect 17500 9172 17552 9178
rect 17184 9132 17264 9160
rect 17132 9114 17184 9120
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 16705 8188 17013 8197
rect 16705 8186 16711 8188
rect 16767 8186 16791 8188
rect 16847 8186 16871 8188
rect 16927 8186 16951 8188
rect 17007 8186 17013 8188
rect 16767 8134 16769 8186
rect 16949 8134 16951 8186
rect 16705 8132 16711 8134
rect 16767 8132 16791 8134
rect 16847 8132 16871 8134
rect 16927 8132 16951 8134
rect 17007 8132 17013 8134
rect 16705 8123 17013 8132
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 17144 7886 17172 8230
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16132 7262 16252 7290
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14752 3942 14780 4490
rect 14844 4078 14872 4490
rect 14936 4486 14964 4966
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 15028 3534 15056 4626
rect 15304 4622 15332 5646
rect 15292 4616 15344 4622
rect 15290 4584 15292 4593
rect 15344 4584 15346 4593
rect 15290 4519 15346 4528
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15212 3194 15240 4082
rect 15396 3534 15424 4422
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15764 3398 15792 6734
rect 15856 6254 15884 6938
rect 16132 6934 16160 7142
rect 16224 7002 16252 7262
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6474 16068 6734
rect 15948 6458 16068 6474
rect 16132 6458 16160 6870
rect 15936 6452 16068 6458
rect 15988 6446 16068 6452
rect 16120 6452 16172 6458
rect 15936 6394 15988 6400
rect 16120 6394 16172 6400
rect 16316 6322 16344 7414
rect 16705 7100 17013 7109
rect 16705 7098 16711 7100
rect 16767 7098 16791 7100
rect 16847 7098 16871 7100
rect 16927 7098 16951 7100
rect 17007 7098 17013 7100
rect 16767 7046 16769 7098
rect 16949 7046 16951 7098
rect 16705 7044 16711 7046
rect 16767 7044 16791 7046
rect 16847 7044 16871 7046
rect 16927 7044 16951 7046
rect 17007 7044 17013 7046
rect 16705 7035 17013 7044
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 15936 6316 15988 6322
rect 16212 6316 16264 6322
rect 15988 6276 16212 6304
rect 15936 6258 15988 6264
rect 16212 6258 16264 6264
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15856 5778 15884 6054
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15948 5250 15976 6054
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16408 5370 16436 5510
rect 16500 5370 16528 6666
rect 16960 6322 17172 6338
rect 17236 6322 17264 9132
rect 17500 9114 17552 9120
rect 17696 8786 17724 9318
rect 17696 8758 17740 8786
rect 17365 8732 17673 8741
rect 17365 8730 17371 8732
rect 17427 8730 17451 8732
rect 17507 8730 17531 8732
rect 17587 8730 17611 8732
rect 17667 8730 17673 8732
rect 17427 8678 17429 8730
rect 17609 8678 17611 8730
rect 17365 8676 17371 8678
rect 17427 8676 17451 8678
rect 17507 8676 17531 8678
rect 17587 8676 17611 8678
rect 17667 8676 17673 8678
rect 17365 8667 17673 8676
rect 17712 8650 17740 8758
rect 17696 8622 17740 8650
rect 17696 7818 17724 8622
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 17365 7644 17673 7653
rect 17365 7642 17371 7644
rect 17427 7642 17451 7644
rect 17507 7642 17531 7644
rect 17587 7642 17611 7644
rect 17667 7642 17673 7644
rect 17427 7590 17429 7642
rect 17609 7590 17611 7642
rect 17365 7588 17371 7590
rect 17427 7588 17451 7590
rect 17507 7588 17531 7590
rect 17587 7588 17611 7590
rect 17667 7588 17673 7590
rect 17365 7579 17673 7588
rect 17788 7018 17816 9540
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17880 8838 17908 9386
rect 18064 8974 18092 9862
rect 18156 9586 18184 9930
rect 18248 9722 18276 11494
rect 18340 11218 18368 11630
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18340 10810 18368 11154
rect 18432 11150 18460 11766
rect 20718 11727 20774 11736
rect 20812 11756 20864 11762
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 11150 19472 11494
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18340 10266 18368 10746
rect 18432 10674 18460 10950
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18340 9466 18368 10202
rect 18524 10198 18552 11086
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18616 10266 18644 10474
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 18708 9654 18736 11018
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10674 18828 10950
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18340 9438 18460 9466
rect 18432 9382 18460 9438
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17880 7886 17908 8774
rect 18156 8498 18184 8774
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 18064 8090 18092 8298
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18248 8022 18276 8910
rect 18340 8498 18368 9318
rect 18432 9178 18460 9318
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18524 8566 18552 8910
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7750 17908 7822
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17880 7410 17908 7686
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17972 7206 18000 7686
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17788 6990 17908 7018
rect 17880 6882 17908 6990
rect 17776 6860 17828 6866
rect 17880 6854 18000 6882
rect 17776 6802 17828 6808
rect 17365 6556 17673 6565
rect 17365 6554 17371 6556
rect 17427 6554 17451 6556
rect 17507 6554 17531 6556
rect 17587 6554 17611 6556
rect 17667 6554 17673 6556
rect 17427 6502 17429 6554
rect 17609 6502 17611 6554
rect 17365 6500 17371 6502
rect 17427 6500 17451 6502
rect 17507 6500 17531 6502
rect 17587 6500 17611 6502
rect 17667 6500 17673 6502
rect 17365 6491 17673 6500
rect 16948 6316 17172 6322
rect 17000 6310 17172 6316
rect 16948 6258 17000 6264
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 15856 5222 15976 5250
rect 15856 5166 15884 5222
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15856 4146 15884 5102
rect 15948 4554 15976 5102
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15948 4146 15976 4490
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 16224 4078 16252 5034
rect 16500 4282 16528 5306
rect 16592 5166 16620 6054
rect 16705 6012 17013 6021
rect 16705 6010 16711 6012
rect 16767 6010 16791 6012
rect 16847 6010 16871 6012
rect 16927 6010 16951 6012
rect 17007 6010 17013 6012
rect 16767 5958 16769 6010
rect 16949 5958 16951 6010
rect 16705 5956 16711 5958
rect 16767 5956 16791 5958
rect 16847 5956 16871 5958
rect 16927 5956 16951 5958
rect 17007 5956 17013 5958
rect 16705 5947 17013 5956
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16684 5030 16712 5510
rect 17052 5098 17080 6190
rect 17144 5914 17172 6310
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17144 5302 17172 5850
rect 17236 5642 17264 6258
rect 17788 5778 17816 6802
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17880 6458 17908 6666
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17972 6338 18000 6854
rect 18156 6798 18184 7958
rect 18340 7546 18368 8230
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18432 7818 18460 8026
rect 18420 7812 18472 7818
rect 18472 7772 18552 7800
rect 18420 7754 18472 7760
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18524 7478 18552 7772
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 17880 6310 18000 6338
rect 18144 6316 18196 6322
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17236 5370 17264 5578
rect 17365 5468 17673 5477
rect 17365 5466 17371 5468
rect 17427 5466 17451 5468
rect 17507 5466 17531 5468
rect 17587 5466 17611 5468
rect 17667 5466 17673 5468
rect 17427 5414 17429 5466
rect 17609 5414 17611 5466
rect 17365 5412 17371 5414
rect 17427 5412 17451 5414
rect 17507 5412 17531 5414
rect 17587 5412 17611 5414
rect 17667 5412 17673 5414
rect 17365 5403 17673 5412
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 5296 17184 5302
rect 17130 5264 17132 5273
rect 17184 5264 17186 5273
rect 17130 5199 17186 5208
rect 17040 5092 17092 5098
rect 17040 5034 17092 5040
rect 17236 5030 17264 5306
rect 17406 5264 17462 5273
rect 17406 5199 17408 5208
rect 17460 5199 17462 5208
rect 17408 5170 17460 5176
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 16592 4622 16620 4966
rect 16705 4924 17013 4933
rect 16705 4922 16711 4924
rect 16767 4922 16791 4924
rect 16847 4922 16871 4924
rect 16927 4922 16951 4924
rect 17007 4922 17013 4924
rect 16767 4870 16769 4922
rect 16949 4870 16951 4922
rect 16705 4868 16711 4870
rect 16767 4868 16791 4870
rect 16847 4868 16871 4870
rect 16927 4868 16951 4870
rect 17007 4868 17013 4870
rect 16705 4859 17013 4868
rect 17420 4622 17448 5170
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16500 3398 16528 4218
rect 16868 4146 16896 4422
rect 17365 4380 17673 4389
rect 17365 4378 17371 4380
rect 17427 4378 17451 4380
rect 17507 4378 17531 4380
rect 17587 4378 17611 4380
rect 17667 4378 17673 4380
rect 17427 4326 17429 4378
rect 17609 4326 17611 4378
rect 17365 4324 17371 4326
rect 17427 4324 17451 4326
rect 17507 4324 17531 4326
rect 17587 4324 17611 4326
rect 17667 4324 17673 4326
rect 17365 4315 17673 4324
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17144 4146 17172 4218
rect 17788 4146 17816 5714
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16705 3836 17013 3845
rect 16705 3834 16711 3836
rect 16767 3834 16791 3836
rect 16847 3834 16871 3836
rect 16927 3834 16951 3836
rect 17007 3834 17013 3836
rect 16767 3782 16769 3834
rect 16949 3782 16951 3834
rect 16705 3780 16711 3782
rect 16767 3780 16791 3782
rect 16847 3780 16871 3782
rect 16927 3780 16951 3782
rect 17007 3780 17013 3782
rect 16705 3771 17013 3780
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 14476 2746 14688 2774
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 14476 2514 14504 2746
rect 16316 2650 16344 2994
rect 17052 2990 17080 3878
rect 17788 3670 17816 4082
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 16705 2748 17013 2757
rect 16705 2746 16711 2748
rect 16767 2746 16791 2748
rect 16847 2746 16871 2748
rect 16927 2746 16951 2748
rect 17007 2746 17013 2748
rect 16767 2694 16769 2746
rect 16949 2694 16951 2746
rect 16705 2692 16711 2694
rect 16767 2692 16791 2694
rect 16847 2692 16871 2694
rect 16927 2692 16951 2694
rect 17007 2692 17013 2694
rect 16705 2683 17013 2692
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 17144 2582 17172 3470
rect 17365 3292 17673 3301
rect 17365 3290 17371 3292
rect 17427 3290 17451 3292
rect 17507 3290 17531 3292
rect 17587 3290 17611 3292
rect 17667 3290 17673 3292
rect 17427 3238 17429 3290
rect 17609 3238 17611 3290
rect 17365 3236 17371 3238
rect 17427 3236 17451 3238
rect 17507 3236 17531 3238
rect 17587 3236 17611 3238
rect 17667 3236 17673 3238
rect 17365 3227 17673 3236
rect 17788 2990 17816 3606
rect 17880 3194 17908 6310
rect 18144 6258 18196 6264
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17972 5710 18000 6122
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18064 5302 18092 5510
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17972 4214 18000 4966
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 18156 3534 18184 6258
rect 18248 3738 18276 7142
rect 18432 7002 18460 7414
rect 18524 7206 18552 7414
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18616 5914 18644 9590
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18708 8974 18736 9386
rect 18892 9382 18920 9522
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18786 9072 18842 9081
rect 18786 9007 18842 9016
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18800 8498 18828 9007
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18984 7818 19012 10610
rect 19076 10062 19104 10610
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19076 8974 19104 9998
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19168 8906 19196 9522
rect 19352 9178 19380 9522
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 19168 7546 19196 8298
rect 19352 7954 19380 8774
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19076 6798 19104 7210
rect 19352 7018 19380 7278
rect 19260 7002 19380 7018
rect 19248 6996 19380 7002
rect 19300 6990 19380 6996
rect 19248 6938 19300 6944
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19076 6254 19104 6734
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 6322 19288 6598
rect 19352 6458 19380 6990
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19338 6216 19394 6225
rect 19338 6151 19340 6160
rect 19392 6151 19394 6160
rect 19340 6122 19392 6128
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 18156 3126 18184 3334
rect 18616 3126 18644 5850
rect 19444 5302 19472 10542
rect 19720 10470 19748 11154
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 20732 10418 20760 11727
rect 20812 11698 20864 11704
rect 20824 11506 20852 11698
rect 21008 11694 21036 12406
rect 21192 12102 21220 12406
rect 21284 12288 21312 12718
rect 21364 12300 21416 12306
rect 21284 12260 21364 12288
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20904 11552 20956 11558
rect 20824 11500 20904 11506
rect 20824 11494 20956 11500
rect 20824 11478 20944 11494
rect 20824 11354 20852 11478
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 21008 10674 21036 11630
rect 21192 11286 21220 11698
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21284 11082 21312 12260
rect 21364 12242 21416 12248
rect 21560 11898 21588 12718
rect 22020 12102 22048 12718
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22296 12170 22324 12582
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21376 11014 21404 11698
rect 21468 11642 21496 11834
rect 21928 11830 21956 12038
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 22020 11778 22048 12038
rect 22192 11824 22244 11830
rect 22020 11772 22192 11778
rect 22020 11766 22244 11772
rect 22020 11762 22232 11766
rect 22388 11762 22416 13126
rect 23124 12986 23152 13194
rect 23667 13084 23975 13093
rect 23667 13082 23673 13084
rect 23729 13082 23753 13084
rect 23809 13082 23833 13084
rect 23889 13082 23913 13084
rect 23969 13082 23975 13084
rect 23729 13030 23731 13082
rect 23911 13030 23913 13082
rect 23667 13028 23673 13030
rect 23729 13028 23753 13030
rect 23809 13028 23833 13030
rect 23889 13028 23913 13030
rect 23969 13028 23975 13030
rect 23667 13019 23975 13028
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23007 12540 23315 12549
rect 23007 12538 23013 12540
rect 23069 12538 23093 12540
rect 23149 12538 23173 12540
rect 23229 12538 23253 12540
rect 23309 12538 23315 12540
rect 23069 12486 23071 12538
rect 23251 12486 23253 12538
rect 23007 12484 23013 12486
rect 23069 12484 23093 12486
rect 23149 12484 23173 12486
rect 23229 12484 23253 12486
rect 23309 12484 23315 12486
rect 23007 12475 23315 12484
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22480 11762 22508 12242
rect 23667 11996 23975 12005
rect 23667 11994 23673 11996
rect 23729 11994 23753 11996
rect 23809 11994 23833 11996
rect 23889 11994 23913 11996
rect 23969 11994 23975 11996
rect 23729 11942 23731 11994
rect 23911 11942 23913 11994
rect 23667 11940 23673 11942
rect 23729 11940 23753 11942
rect 23809 11940 23833 11942
rect 23889 11940 23913 11942
rect 23969 11940 23975 11942
rect 23667 11931 23975 11940
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23110 11792 23166 11801
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 22008 11756 22232 11762
rect 22060 11750 22232 11756
rect 22376 11756 22428 11762
rect 22008 11698 22060 11704
rect 22296 11716 22376 11744
rect 21468 11614 21588 11642
rect 21560 11608 21588 11614
rect 21640 11620 21692 11626
rect 21560 11580 21640 11608
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21468 11150 21496 11494
rect 21560 11150 21588 11580
rect 21640 11562 21692 11568
rect 21836 11558 21864 11698
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 21836 11150 21864 11494
rect 22020 11218 22048 11494
rect 22296 11354 22324 11716
rect 22376 11698 22428 11704
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22928 11756 22980 11762
rect 23110 11727 23112 11736
rect 22928 11698 22980 11704
rect 23164 11727 23166 11736
rect 23112 11698 23164 11704
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 10674 21404 10950
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21088 10464 21140 10470
rect 19720 10062 19748 10406
rect 20732 10390 20852 10418
rect 21088 10406 21140 10412
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20640 9654 20668 9998
rect 20732 9654 20760 10134
rect 20824 10130 20852 10390
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20640 9466 20668 9590
rect 20640 9450 20760 9466
rect 20640 9444 20772 9450
rect 20640 9438 20720 9444
rect 20720 9386 20772 9392
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19536 7342 19564 7958
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19536 6322 19564 6394
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19536 5846 19564 6258
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19444 4758 19472 5238
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19432 4616 19484 4622
rect 19536 4604 19564 5238
rect 19628 5030 19656 9318
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 19720 8090 19748 9046
rect 20824 9042 20852 10066
rect 20916 9364 20944 10202
rect 21100 10130 21128 10406
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 21008 9586 21036 9930
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21376 9586 21404 9862
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21468 9518 21496 10610
rect 21560 9586 21588 11086
rect 22020 10674 22048 11154
rect 22204 10810 22232 11154
rect 22940 11150 22968 11698
rect 23007 11452 23315 11461
rect 23007 11450 23013 11452
rect 23069 11450 23093 11452
rect 23149 11450 23173 11452
rect 23229 11450 23253 11452
rect 23309 11450 23315 11452
rect 23069 11398 23071 11450
rect 23251 11398 23253 11450
rect 23007 11396 23013 11398
rect 23069 11396 23093 11398
rect 23149 11396 23173 11398
rect 23229 11396 23253 11398
rect 23309 11396 23315 11398
rect 23007 11387 23315 11396
rect 23492 11218 23520 11834
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21836 9586 21864 10202
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22112 9586 22140 9658
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21560 9382 21588 9522
rect 20996 9376 21048 9382
rect 20916 9336 20996 9364
rect 20996 9318 21048 9324
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21008 9178 21036 9318
rect 22112 9178 22140 9522
rect 22296 9382 22324 10610
rect 22940 10266 22968 11086
rect 23492 10606 23520 11154
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23007 10364 23315 10373
rect 23007 10362 23013 10364
rect 23069 10362 23093 10364
rect 23149 10362 23173 10364
rect 23229 10362 23253 10364
rect 23309 10362 23315 10364
rect 23069 10310 23071 10362
rect 23251 10310 23253 10362
rect 23007 10308 23013 10310
rect 23069 10308 23093 10310
rect 23149 10308 23173 10310
rect 23229 10308 23253 10310
rect 23309 10308 23315 10310
rect 23007 10299 23315 10308
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 22376 9988 22428 9994
rect 22376 9930 22428 9936
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22388 9178 22416 9930
rect 23308 9926 23336 9998
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 22572 9586 22600 9862
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 23308 9450 23336 9862
rect 23400 9722 23428 9998
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23400 9602 23428 9658
rect 23400 9574 23520 9602
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 22468 9444 22520 9450
rect 22468 9386 22520 9392
rect 23296 9444 23348 9450
rect 23296 9386 23348 9392
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22480 9110 22508 9386
rect 23007 9276 23315 9285
rect 23007 9274 23013 9276
rect 23069 9274 23093 9276
rect 23149 9274 23173 9276
rect 23229 9274 23253 9276
rect 23309 9274 23315 9276
rect 23069 9222 23071 9274
rect 23251 9222 23253 9274
rect 23007 9220 23013 9222
rect 23069 9220 23093 9222
rect 23149 9220 23173 9222
rect 23229 9220 23253 9222
rect 23309 9220 23315 9222
rect 23007 9211 23315 9220
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8634 20300 8910
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20824 8566 20852 8978
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 22480 8362 22508 9046
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22572 8498 22600 8910
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22664 8634 22692 8842
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 23400 8498 23428 9454
rect 23492 9382 23520 9574
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23584 8566 23612 11222
rect 23952 11132 23980 11494
rect 24044 11354 24072 11630
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24032 11144 24084 11150
rect 23952 11104 24032 11132
rect 24032 11086 24084 11092
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 23667 10908 23975 10917
rect 23667 10906 23673 10908
rect 23729 10906 23753 10908
rect 23809 10906 23833 10908
rect 23889 10906 23913 10908
rect 23969 10906 23975 10908
rect 23729 10854 23731 10906
rect 23911 10854 23913 10906
rect 23667 10852 23673 10854
rect 23729 10852 23753 10854
rect 23809 10852 23833 10854
rect 23889 10852 23913 10854
rect 23969 10852 23975 10854
rect 23667 10843 23975 10852
rect 24136 10810 24164 11018
rect 24228 11014 24256 11086
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24124 10804 24176 10810
rect 24124 10746 24176 10752
rect 24228 10674 24256 10950
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 23676 9994 23704 10610
rect 23860 10198 23888 10610
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23667 9820 23975 9829
rect 23667 9818 23673 9820
rect 23729 9818 23753 9820
rect 23809 9818 23833 9820
rect 23889 9818 23913 9820
rect 23969 9818 23975 9820
rect 23729 9766 23731 9818
rect 23911 9766 23913 9818
rect 23667 9764 23673 9766
rect 23729 9764 23753 9766
rect 23809 9764 23833 9766
rect 23889 9764 23913 9766
rect 23969 9764 23975 9766
rect 23667 9755 23975 9764
rect 24136 9654 24164 10406
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 23667 8732 23975 8741
rect 23667 8730 23673 8732
rect 23729 8730 23753 8732
rect 23809 8730 23833 8732
rect 23889 8730 23913 8732
rect 23969 8730 23975 8732
rect 23729 8678 23731 8730
rect 23911 8678 23913 8730
rect 23667 8676 23673 8678
rect 23729 8676 23753 8678
rect 23809 8676 23833 8678
rect 23889 8676 23913 8678
rect 23969 8676 23975 8678
rect 23667 8667 23975 8676
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 23007 8188 23315 8197
rect 23007 8186 23013 8188
rect 23069 8186 23093 8188
rect 23149 8186 23173 8188
rect 23229 8186 23253 8188
rect 23309 8186 23315 8188
rect 23069 8134 23071 8186
rect 23251 8134 23253 8186
rect 23007 8132 23013 8134
rect 23069 8132 23093 8134
rect 23149 8132 23173 8134
rect 23229 8132 23253 8134
rect 23309 8132 23315 8134
rect 23007 8123 23315 8132
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19720 6458 19748 6734
rect 19812 6662 19840 7414
rect 21468 7410 21496 7686
rect 22664 7546 22692 7822
rect 23667 7644 23975 7653
rect 23667 7642 23673 7644
rect 23729 7642 23753 7644
rect 23809 7642 23833 7644
rect 23889 7642 23913 7644
rect 23969 7642 23975 7644
rect 23729 7590 23731 7642
rect 23911 7590 23913 7642
rect 23667 7588 23673 7590
rect 23729 7588 23753 7590
rect 23809 7588 23833 7590
rect 23889 7588 23913 7590
rect 23969 7588 23975 7590
rect 23667 7579 23975 7588
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 20628 7336 20680 7342
rect 20548 7296 20628 7324
rect 20548 7002 20576 7296
rect 20628 7278 20680 7284
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20824 7002 20852 7278
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19706 6352 19762 6361
rect 19706 6287 19708 6296
rect 19760 6287 19762 6296
rect 19708 6258 19760 6264
rect 19812 6118 19840 6598
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19996 6118 20024 6326
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 19708 6112 19760 6118
rect 19706 6080 19708 6089
rect 19800 6112 19852 6118
rect 19760 6080 19762 6089
rect 19800 6054 19852 6060
rect 19984 6112 20036 6118
rect 20036 6072 20116 6100
rect 19984 6054 20036 6060
rect 19706 6015 19762 6024
rect 19984 5296 20036 5302
rect 19984 5238 20036 5244
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19628 4690 19656 4966
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 19484 4576 19564 4604
rect 19432 4558 19484 4564
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 19260 4078 19288 4422
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19352 3534 19380 4150
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18892 2990 18920 3470
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 19444 2922 19472 4558
rect 19996 4554 20024 5238
rect 20088 5114 20116 6072
rect 20180 5681 20208 6258
rect 20352 6248 20404 6254
rect 20350 6216 20352 6225
rect 20404 6216 20406 6225
rect 20350 6151 20406 6160
rect 20260 5704 20312 5710
rect 20166 5672 20222 5681
rect 20260 5646 20312 5652
rect 20166 5607 20222 5616
rect 20272 5370 20300 5646
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20456 5166 20484 6258
rect 20548 6089 20576 6938
rect 20824 6361 20852 6938
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 20810 6352 20866 6361
rect 20810 6287 20866 6296
rect 20996 6316 21048 6322
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20534 6080 20590 6089
rect 20534 6015 20590 6024
rect 20640 5914 20668 6190
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20824 5642 20852 6287
rect 20996 6258 21048 6264
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 21008 5370 21036 6258
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 20444 5160 20496 5166
rect 20088 5086 20300 5114
rect 20444 5102 20496 5108
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19996 4282 20024 4490
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 20088 4078 20116 4966
rect 20168 4752 20220 4758
rect 20168 4694 20220 4700
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19628 3534 19656 3946
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19904 3058 19932 3334
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 20180 2990 20208 4694
rect 20272 4690 20300 5086
rect 20456 4690 20484 5102
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20824 4690 20852 4966
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20272 4486 20300 4626
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20260 4140 20312 4146
rect 20456 4128 20484 4626
rect 20824 4282 20852 4626
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20536 4140 20588 4146
rect 20456 4100 20536 4128
rect 20260 4082 20312 4088
rect 20536 4082 20588 4088
rect 20272 3194 20300 4082
rect 20824 3738 20852 4218
rect 21008 4078 21036 4422
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20444 3460 20496 3466
rect 20444 3402 20496 3408
rect 20456 3194 20484 3402
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20824 3126 20852 3674
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 21192 3058 21220 6734
rect 21284 6322 21312 7142
rect 21928 6866 21956 7346
rect 22572 6866 22600 7414
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21928 6254 21956 6802
rect 22664 6440 22692 7482
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 23007 7100 23315 7109
rect 23007 7098 23013 7100
rect 23069 7098 23093 7100
rect 23149 7098 23173 7100
rect 23229 7098 23253 7100
rect 23309 7098 23315 7100
rect 23069 7046 23071 7098
rect 23251 7046 23253 7098
rect 23007 7044 23013 7046
rect 23069 7044 23093 7046
rect 23149 7044 23173 7046
rect 23229 7044 23253 7046
rect 23309 7044 23315 7046
rect 23007 7035 23315 7044
rect 24044 6798 24072 7414
rect 24320 7410 24348 15302
rect 25056 13530 25084 18226
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25700 16794 25728 17138
rect 25870 17096 25926 17105
rect 25870 17031 25872 17040
rect 25924 17031 25926 17040
rect 25872 17002 25924 17008
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25792 13025 25820 13262
rect 25778 13016 25834 13025
rect 25778 12951 25834 12960
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24688 12238 24716 12786
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24504 11830 24532 12038
rect 24492 11824 24544 11830
rect 24492 11766 24544 11772
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24504 10266 24532 10610
rect 24596 10606 24624 11698
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24688 10130 24716 12174
rect 24952 11620 25004 11626
rect 24952 11562 25004 11568
rect 24964 10674 24992 11562
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25700 11218 25728 11494
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 24780 10266 24808 10610
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24504 9994 24532 10066
rect 24492 9988 24544 9994
rect 24492 9930 24544 9936
rect 24688 8974 24716 10066
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 24872 9518 24900 9998
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 25148 9382 25176 9998
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25424 9654 25452 9862
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 24412 8566 24440 8774
rect 24400 8560 24452 8566
rect 24400 8502 24452 8508
rect 24688 7478 24716 8910
rect 25148 8634 25176 9318
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25872 8356 25924 8362
rect 25872 8298 25924 8304
rect 25884 8265 25912 8298
rect 25870 8256 25926 8265
rect 25870 8191 25926 8200
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 22572 6412 22692 6440
rect 22572 6322 22600 6412
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21652 4622 21680 5850
rect 21928 5778 21956 6190
rect 22388 6118 22416 6258
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22284 6112 22336 6118
rect 22376 6112 22428 6118
rect 22284 6054 22336 6060
rect 22374 6080 22376 6089
rect 22428 6080 22430 6089
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 22020 5642 22048 6054
rect 22296 5710 22324 6054
rect 22374 6015 22430 6024
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22284 5704 22336 5710
rect 22572 5681 22600 5714
rect 22284 5646 22336 5652
rect 22558 5672 22614 5681
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 22008 5636 22060 5642
rect 22008 5578 22060 5584
rect 21744 4690 21772 5578
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 4146 21680 4558
rect 22020 4554 22048 5170
rect 22008 4548 22060 4554
rect 22008 4490 22060 4496
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 22296 4078 22324 5646
rect 22558 5607 22614 5616
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22388 4486 22416 5510
rect 22572 5234 22600 5607
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22480 4214 22508 4422
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 22376 4140 22428 4146
rect 22572 4128 22600 5170
rect 22664 5098 22692 6258
rect 22756 5710 22784 6258
rect 22940 5914 22968 6258
rect 23007 6012 23315 6021
rect 23007 6010 23013 6012
rect 23069 6010 23093 6012
rect 23149 6010 23173 6012
rect 23229 6010 23253 6012
rect 23309 6010 23315 6012
rect 23069 5958 23071 6010
rect 23251 5958 23253 6010
rect 23007 5956 23013 5958
rect 23069 5956 23093 5958
rect 23149 5956 23173 5958
rect 23229 5956 23253 5958
rect 23309 5956 23315 5958
rect 23007 5947 23315 5956
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22756 5370 22784 5646
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22940 5234 22968 5850
rect 23584 5642 23612 6598
rect 23667 6556 23975 6565
rect 23667 6554 23673 6556
rect 23729 6554 23753 6556
rect 23809 6554 23833 6556
rect 23889 6554 23913 6556
rect 23969 6554 23975 6556
rect 23729 6502 23731 6554
rect 23911 6502 23913 6554
rect 23667 6500 23673 6502
rect 23729 6500 23753 6502
rect 23809 6500 23833 6502
rect 23889 6500 23913 6502
rect 23969 6500 23975 6502
rect 23667 6491 23975 6500
rect 24136 6390 24164 6598
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 23572 5636 23624 5642
rect 23572 5578 23624 5584
rect 23667 5468 23975 5477
rect 23667 5466 23673 5468
rect 23729 5466 23753 5468
rect 23809 5466 23833 5468
rect 23889 5466 23913 5468
rect 23969 5466 23975 5468
rect 23729 5414 23731 5466
rect 23911 5414 23913 5466
rect 23667 5412 23673 5414
rect 23729 5412 23753 5414
rect 23809 5412 23833 5414
rect 23889 5412 23913 5414
rect 23969 5412 23975 5414
rect 23667 5403 23975 5412
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22652 5092 22704 5098
rect 22652 5034 22704 5040
rect 22848 4978 22876 5170
rect 22848 4950 22968 4978
rect 22940 4214 22968 4950
rect 23007 4924 23315 4933
rect 23007 4922 23013 4924
rect 23069 4922 23093 4924
rect 23149 4922 23173 4924
rect 23229 4922 23253 4924
rect 23309 4922 23315 4924
rect 23069 4870 23071 4922
rect 23251 4870 23253 4922
rect 23007 4868 23013 4870
rect 23069 4868 23093 4870
rect 23149 4868 23173 4870
rect 23229 4868 23253 4870
rect 23309 4868 23315 4870
rect 23007 4859 23315 4868
rect 23667 4380 23975 4389
rect 23667 4378 23673 4380
rect 23729 4378 23753 4380
rect 23809 4378 23833 4380
rect 23889 4378 23913 4380
rect 23969 4378 23975 4380
rect 23729 4326 23731 4378
rect 23911 4326 23913 4378
rect 23667 4324 23673 4326
rect 23729 4324 23753 4326
rect 23809 4324 23833 4326
rect 23889 4324 23913 4326
rect 23969 4324 23975 4326
rect 23667 4315 23975 4324
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 22652 4140 22704 4146
rect 22572 4100 22652 4128
rect 22376 4082 22428 4088
rect 22652 4082 22704 4088
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22388 3738 22416 4082
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22664 3602 22692 3878
rect 23007 3836 23315 3845
rect 23007 3834 23013 3836
rect 23069 3834 23093 3836
rect 23149 3834 23173 3836
rect 23229 3834 23253 3836
rect 23309 3834 23315 3836
rect 23069 3782 23071 3834
rect 23251 3782 23253 3834
rect 23007 3780 23013 3782
rect 23069 3780 23093 3782
rect 23149 3780 23173 3782
rect 23229 3780 23253 3782
rect 23309 3780 23315 3782
rect 23007 3771 23315 3780
rect 24320 3738 24348 7346
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 25792 4185 25820 4558
rect 25778 4176 25834 4185
rect 25778 4111 25834 4120
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 21928 3194 21956 3402
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 23007 2748 23315 2757
rect 23007 2746 23013 2748
rect 23069 2746 23093 2748
rect 23149 2746 23173 2748
rect 23229 2746 23253 2748
rect 23309 2746 23315 2748
rect 23069 2694 23071 2746
rect 23251 2694 23253 2746
rect 23007 2692 23013 2694
rect 23069 2692 23093 2694
rect 23149 2692 23173 2694
rect 23229 2692 23253 2694
rect 23309 2692 23315 2694
rect 23007 2683 23315 2692
rect 23584 2650 23612 3470
rect 23667 3292 23975 3301
rect 23667 3290 23673 3292
rect 23729 3290 23753 3292
rect 23809 3290 23833 3292
rect 23889 3290 23913 3292
rect 23969 3290 23975 3292
rect 23729 3238 23731 3290
rect 23911 3238 23913 3290
rect 23667 3236 23673 3238
rect 23729 3236 23753 3238
rect 23809 3236 23833 3238
rect 23889 3236 23913 3238
rect 23969 3236 23975 3238
rect 23667 3227 23975 3236
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 15488 800 15516 2382
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 17365 2204 17673 2213
rect 17365 2202 17371 2204
rect 17427 2202 17451 2204
rect 17507 2202 17531 2204
rect 17587 2202 17611 2204
rect 17667 2202 17673 2204
rect 17427 2150 17429 2202
rect 17609 2150 17611 2202
rect 17365 2148 17371 2150
rect 17427 2148 17451 2150
rect 17507 2148 17531 2150
rect 17587 2148 17611 2150
rect 17667 2148 17673 2150
rect 17365 2139 17673 2148
rect 19996 800 20024 2246
rect 23667 2204 23975 2213
rect 23667 2202 23673 2204
rect 23729 2202 23753 2204
rect 23809 2202 23833 2204
rect 23889 2202 23913 2204
rect 23969 2202 23975 2204
rect 23729 2150 23731 2202
rect 23911 2150 23913 2202
rect 23667 2148 23673 2150
rect 23729 2148 23753 2150
rect 23809 2148 23833 2150
rect 23889 2148 23913 2150
rect 23969 2148 23975 2150
rect 23667 2139 23975 2148
rect 24044 1306 24072 2382
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 23860 1278 24072 1306
rect 23860 800 23888 1278
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
rect 19982 0 20038 800
rect 23846 0 23902 800
rect 24780 105 24808 2246
rect 24766 96 24822 105
rect 24766 31 24822 40
<< via2 >>
rect 1398 29280 1454 29336
rect 4767 27226 4823 27228
rect 4847 27226 4903 27228
rect 4927 27226 4983 27228
rect 5007 27226 5063 27228
rect 4767 27174 4813 27226
rect 4813 27174 4823 27226
rect 4847 27174 4877 27226
rect 4877 27174 4889 27226
rect 4889 27174 4903 27226
rect 4927 27174 4941 27226
rect 4941 27174 4953 27226
rect 4953 27174 4983 27226
rect 5007 27174 5017 27226
rect 5017 27174 5063 27226
rect 4767 27172 4823 27174
rect 4847 27172 4903 27174
rect 4927 27172 4983 27174
rect 5007 27172 5063 27174
rect 11069 27226 11125 27228
rect 11149 27226 11205 27228
rect 11229 27226 11285 27228
rect 11309 27226 11365 27228
rect 11069 27174 11115 27226
rect 11115 27174 11125 27226
rect 11149 27174 11179 27226
rect 11179 27174 11191 27226
rect 11191 27174 11205 27226
rect 11229 27174 11243 27226
rect 11243 27174 11255 27226
rect 11255 27174 11285 27226
rect 11309 27174 11319 27226
rect 11319 27174 11365 27226
rect 11069 27172 11125 27174
rect 11149 27172 11205 27174
rect 11229 27172 11285 27174
rect 11309 27172 11365 27174
rect 938 21120 994 21176
rect 1582 20440 1638 20496
rect 4107 26682 4163 26684
rect 4187 26682 4243 26684
rect 4267 26682 4323 26684
rect 4347 26682 4403 26684
rect 4107 26630 4153 26682
rect 4153 26630 4163 26682
rect 4187 26630 4217 26682
rect 4217 26630 4229 26682
rect 4229 26630 4243 26682
rect 4267 26630 4281 26682
rect 4281 26630 4293 26682
rect 4293 26630 4323 26682
rect 4347 26630 4357 26682
rect 4357 26630 4403 26682
rect 4107 26628 4163 26630
rect 4187 26628 4243 26630
rect 4267 26628 4323 26630
rect 4347 26628 4403 26630
rect 10409 26682 10465 26684
rect 10489 26682 10545 26684
rect 10569 26682 10625 26684
rect 10649 26682 10705 26684
rect 10409 26630 10455 26682
rect 10455 26630 10465 26682
rect 10489 26630 10519 26682
rect 10519 26630 10531 26682
rect 10531 26630 10545 26682
rect 10569 26630 10583 26682
rect 10583 26630 10595 26682
rect 10595 26630 10625 26682
rect 10649 26630 10659 26682
rect 10659 26630 10705 26682
rect 10409 26628 10465 26630
rect 10489 26628 10545 26630
rect 10569 26628 10625 26630
rect 10649 26628 10705 26630
rect 4767 26138 4823 26140
rect 4847 26138 4903 26140
rect 4927 26138 4983 26140
rect 5007 26138 5063 26140
rect 4767 26086 4813 26138
rect 4813 26086 4823 26138
rect 4847 26086 4877 26138
rect 4877 26086 4889 26138
rect 4889 26086 4903 26138
rect 4927 26086 4941 26138
rect 4941 26086 4953 26138
rect 4953 26086 4983 26138
rect 5007 26086 5017 26138
rect 5017 26086 5063 26138
rect 4767 26084 4823 26086
rect 4847 26084 4903 26086
rect 4927 26084 4983 26086
rect 5007 26084 5063 26086
rect 4107 25594 4163 25596
rect 4187 25594 4243 25596
rect 4267 25594 4323 25596
rect 4347 25594 4403 25596
rect 4107 25542 4153 25594
rect 4153 25542 4163 25594
rect 4187 25542 4217 25594
rect 4217 25542 4229 25594
rect 4229 25542 4243 25594
rect 4267 25542 4281 25594
rect 4281 25542 4293 25594
rect 4293 25542 4323 25594
rect 4347 25542 4357 25594
rect 4357 25542 4403 25594
rect 4107 25540 4163 25542
rect 4187 25540 4243 25542
rect 4267 25540 4323 25542
rect 4347 25540 4403 25542
rect 3238 25200 3294 25256
rect 2594 19760 2650 19816
rect 938 16360 994 16416
rect 4767 25050 4823 25052
rect 4847 25050 4903 25052
rect 4927 25050 4983 25052
rect 5007 25050 5063 25052
rect 4767 24998 4813 25050
rect 4813 24998 4823 25050
rect 4847 24998 4877 25050
rect 4877 24998 4889 25050
rect 4889 24998 4903 25050
rect 4927 24998 4941 25050
rect 4941 24998 4953 25050
rect 4953 24998 4983 25050
rect 5007 24998 5017 25050
rect 5017 24998 5063 25050
rect 4767 24996 4823 24998
rect 4847 24996 4903 24998
rect 4927 24996 4983 24998
rect 5007 24996 5063 24998
rect 4107 24506 4163 24508
rect 4187 24506 4243 24508
rect 4267 24506 4323 24508
rect 4347 24506 4403 24508
rect 4107 24454 4153 24506
rect 4153 24454 4163 24506
rect 4187 24454 4217 24506
rect 4217 24454 4229 24506
rect 4229 24454 4243 24506
rect 4267 24454 4281 24506
rect 4281 24454 4293 24506
rect 4293 24454 4323 24506
rect 4347 24454 4357 24506
rect 4357 24454 4403 24506
rect 4107 24452 4163 24454
rect 4187 24452 4243 24454
rect 4267 24452 4323 24454
rect 4347 24452 4403 24454
rect 4767 23962 4823 23964
rect 4847 23962 4903 23964
rect 4927 23962 4983 23964
rect 5007 23962 5063 23964
rect 4767 23910 4813 23962
rect 4813 23910 4823 23962
rect 4847 23910 4877 23962
rect 4877 23910 4889 23962
rect 4889 23910 4903 23962
rect 4927 23910 4941 23962
rect 4941 23910 4953 23962
rect 4953 23910 4983 23962
rect 5007 23910 5017 23962
rect 5017 23910 5063 23962
rect 4767 23908 4823 23910
rect 4847 23908 4903 23910
rect 4927 23908 4983 23910
rect 5007 23908 5063 23910
rect 5170 23740 5172 23760
rect 5172 23740 5224 23760
rect 5224 23740 5226 23760
rect 5170 23704 5226 23740
rect 6458 23568 6514 23624
rect 6826 23568 6882 23624
rect 1582 12280 1638 12336
rect 1398 8200 1454 8256
rect 5538 23432 5594 23488
rect 4107 23418 4163 23420
rect 4187 23418 4243 23420
rect 4267 23418 4323 23420
rect 4347 23418 4403 23420
rect 4107 23366 4153 23418
rect 4153 23366 4163 23418
rect 4187 23366 4217 23418
rect 4217 23366 4229 23418
rect 4229 23366 4243 23418
rect 4267 23366 4281 23418
rect 4281 23366 4293 23418
rect 4293 23366 4323 23418
rect 4347 23366 4357 23418
rect 4357 23366 4403 23418
rect 4107 23364 4163 23366
rect 4187 23364 4243 23366
rect 4267 23364 4323 23366
rect 4347 23364 4403 23366
rect 4767 22874 4823 22876
rect 4847 22874 4903 22876
rect 4927 22874 4983 22876
rect 5007 22874 5063 22876
rect 4767 22822 4813 22874
rect 4813 22822 4823 22874
rect 4847 22822 4877 22874
rect 4877 22822 4889 22874
rect 4889 22822 4903 22874
rect 4927 22822 4941 22874
rect 4941 22822 4953 22874
rect 4953 22822 4983 22874
rect 5007 22822 5017 22874
rect 5017 22822 5063 22874
rect 4767 22820 4823 22822
rect 4847 22820 4903 22822
rect 4927 22820 4983 22822
rect 5007 22820 5063 22822
rect 9126 25236 9128 25256
rect 9128 25236 9180 25256
rect 9180 25236 9182 25256
rect 9126 25200 9182 25236
rect 10409 25594 10465 25596
rect 10489 25594 10545 25596
rect 10569 25594 10625 25596
rect 10649 25594 10705 25596
rect 10409 25542 10455 25594
rect 10455 25542 10465 25594
rect 10489 25542 10519 25594
rect 10519 25542 10531 25594
rect 10531 25542 10545 25594
rect 10569 25542 10583 25594
rect 10583 25542 10595 25594
rect 10595 25542 10625 25594
rect 10649 25542 10659 25594
rect 10659 25542 10705 25594
rect 10409 25540 10465 25542
rect 10489 25540 10545 25542
rect 10569 25540 10625 25542
rect 10649 25540 10705 25542
rect 10138 25200 10194 25256
rect 9310 23840 9366 23896
rect 9494 23432 9550 23488
rect 9954 24012 9956 24032
rect 9956 24012 10008 24032
rect 10008 24012 10010 24032
rect 9954 23976 10010 24012
rect 10046 23840 10102 23896
rect 10409 24506 10465 24508
rect 10489 24506 10545 24508
rect 10569 24506 10625 24508
rect 10649 24506 10705 24508
rect 10409 24454 10455 24506
rect 10455 24454 10465 24506
rect 10489 24454 10519 24506
rect 10519 24454 10531 24506
rect 10531 24454 10545 24506
rect 10569 24454 10583 24506
rect 10583 24454 10595 24506
rect 10595 24454 10625 24506
rect 10649 24454 10659 24506
rect 10659 24454 10705 24506
rect 10409 24452 10465 24454
rect 10489 24452 10545 24454
rect 10569 24452 10625 24454
rect 10649 24452 10705 24454
rect 10690 23976 10746 24032
rect 17371 27226 17427 27228
rect 17451 27226 17507 27228
rect 17531 27226 17587 27228
rect 17611 27226 17667 27228
rect 17371 27174 17417 27226
rect 17417 27174 17427 27226
rect 17451 27174 17481 27226
rect 17481 27174 17493 27226
rect 17493 27174 17507 27226
rect 17531 27174 17545 27226
rect 17545 27174 17557 27226
rect 17557 27174 17587 27226
rect 17611 27174 17621 27226
rect 17621 27174 17667 27226
rect 17371 27172 17427 27174
rect 17451 27172 17507 27174
rect 17531 27172 17587 27174
rect 17611 27172 17667 27174
rect 23673 27226 23729 27228
rect 23753 27226 23809 27228
rect 23833 27226 23889 27228
rect 23913 27226 23969 27228
rect 23673 27174 23719 27226
rect 23719 27174 23729 27226
rect 23753 27174 23783 27226
rect 23783 27174 23795 27226
rect 23795 27174 23809 27226
rect 23833 27174 23847 27226
rect 23847 27174 23859 27226
rect 23859 27174 23889 27226
rect 23913 27174 23923 27226
rect 23923 27174 23969 27226
rect 23673 27172 23729 27174
rect 23753 27172 23809 27174
rect 23833 27172 23889 27174
rect 23913 27172 23969 27174
rect 11069 26138 11125 26140
rect 11149 26138 11205 26140
rect 11229 26138 11285 26140
rect 11309 26138 11365 26140
rect 11069 26086 11115 26138
rect 11115 26086 11125 26138
rect 11149 26086 11179 26138
rect 11179 26086 11191 26138
rect 11191 26086 11205 26138
rect 11229 26086 11243 26138
rect 11243 26086 11255 26138
rect 11255 26086 11285 26138
rect 11309 26086 11319 26138
rect 11319 26086 11365 26138
rect 11069 26084 11125 26086
rect 11149 26084 11205 26086
rect 11229 26084 11285 26086
rect 11309 26084 11365 26086
rect 11069 25050 11125 25052
rect 11149 25050 11205 25052
rect 11229 25050 11285 25052
rect 11309 25050 11365 25052
rect 11069 24998 11115 25050
rect 11115 24998 11125 25050
rect 11149 24998 11179 25050
rect 11179 24998 11191 25050
rect 11191 24998 11205 25050
rect 11229 24998 11243 25050
rect 11243 24998 11255 25050
rect 11255 24998 11285 25050
rect 11309 24998 11319 25050
rect 11319 24998 11365 25050
rect 11069 24996 11125 24998
rect 11149 24996 11205 24998
rect 11229 24996 11285 24998
rect 11309 24996 11365 24998
rect 11069 23962 11125 23964
rect 11149 23962 11205 23964
rect 11229 23962 11285 23964
rect 11309 23962 11365 23964
rect 11069 23910 11115 23962
rect 11115 23910 11125 23962
rect 11149 23910 11179 23962
rect 11179 23910 11191 23962
rect 11191 23910 11205 23962
rect 11229 23910 11243 23962
rect 11243 23910 11255 23962
rect 11255 23910 11285 23962
rect 11309 23910 11319 23962
rect 11319 23910 11365 23962
rect 11069 23908 11125 23910
rect 11149 23908 11205 23910
rect 11229 23908 11285 23910
rect 11309 23908 11365 23910
rect 9954 23296 10010 23352
rect 10138 23432 10194 23488
rect 10409 23418 10465 23420
rect 10489 23418 10545 23420
rect 10569 23418 10625 23420
rect 10649 23418 10705 23420
rect 10409 23366 10455 23418
rect 10455 23366 10465 23418
rect 10489 23366 10519 23418
rect 10519 23366 10531 23418
rect 10531 23366 10545 23418
rect 10569 23366 10583 23418
rect 10583 23366 10595 23418
rect 10595 23366 10625 23418
rect 10649 23366 10659 23418
rect 10659 23366 10705 23418
rect 10409 23364 10465 23366
rect 10489 23364 10545 23366
rect 10569 23364 10625 23366
rect 10649 23364 10705 23366
rect 10782 23160 10838 23216
rect 11058 23568 11114 23624
rect 11069 22874 11125 22876
rect 11149 22874 11205 22876
rect 11229 22874 11285 22876
rect 11309 22874 11365 22876
rect 11069 22822 11115 22874
rect 11115 22822 11125 22874
rect 11149 22822 11179 22874
rect 11179 22822 11191 22874
rect 11191 22822 11205 22874
rect 11229 22822 11243 22874
rect 11243 22822 11255 22874
rect 11255 22822 11285 22874
rect 11309 22822 11319 22874
rect 11319 22822 11365 22874
rect 11069 22820 11125 22822
rect 11149 22820 11205 22822
rect 11229 22820 11285 22822
rect 11309 22820 11365 22822
rect 4107 22330 4163 22332
rect 4187 22330 4243 22332
rect 4267 22330 4323 22332
rect 4347 22330 4403 22332
rect 4107 22278 4153 22330
rect 4153 22278 4163 22330
rect 4187 22278 4217 22330
rect 4217 22278 4229 22330
rect 4229 22278 4243 22330
rect 4267 22278 4281 22330
rect 4281 22278 4293 22330
rect 4293 22278 4323 22330
rect 4347 22278 4357 22330
rect 4357 22278 4403 22330
rect 4107 22276 4163 22278
rect 4187 22276 4243 22278
rect 4267 22276 4323 22278
rect 4347 22276 4403 22278
rect 4158 21972 4160 21992
rect 4160 21972 4212 21992
rect 4212 21972 4214 21992
rect 4158 21936 4214 21972
rect 4894 21936 4950 21992
rect 4767 21786 4823 21788
rect 4847 21786 4903 21788
rect 4927 21786 4983 21788
rect 5007 21786 5063 21788
rect 4767 21734 4813 21786
rect 4813 21734 4823 21786
rect 4847 21734 4877 21786
rect 4877 21734 4889 21786
rect 4889 21734 4903 21786
rect 4927 21734 4941 21786
rect 4941 21734 4953 21786
rect 4953 21734 4983 21786
rect 5007 21734 5017 21786
rect 5017 21734 5063 21786
rect 4767 21732 4823 21734
rect 4847 21732 4903 21734
rect 4927 21732 4983 21734
rect 5007 21732 5063 21734
rect 4107 21242 4163 21244
rect 4187 21242 4243 21244
rect 4267 21242 4323 21244
rect 4347 21242 4403 21244
rect 4107 21190 4153 21242
rect 4153 21190 4163 21242
rect 4187 21190 4217 21242
rect 4217 21190 4229 21242
rect 4229 21190 4243 21242
rect 4267 21190 4281 21242
rect 4281 21190 4293 21242
rect 4293 21190 4323 21242
rect 4347 21190 4357 21242
rect 4357 21190 4403 21242
rect 4107 21188 4163 21190
rect 4187 21188 4243 21190
rect 4267 21188 4323 21190
rect 4347 21188 4403 21190
rect 4767 20698 4823 20700
rect 4847 20698 4903 20700
rect 4927 20698 4983 20700
rect 5007 20698 5063 20700
rect 4767 20646 4813 20698
rect 4813 20646 4823 20698
rect 4847 20646 4877 20698
rect 4877 20646 4889 20698
rect 4889 20646 4903 20698
rect 4927 20646 4941 20698
rect 4941 20646 4953 20698
rect 4953 20646 4983 20698
rect 5007 20646 5017 20698
rect 5017 20646 5063 20698
rect 4767 20644 4823 20646
rect 4847 20644 4903 20646
rect 4927 20644 4983 20646
rect 5007 20644 5063 20646
rect 4107 20154 4163 20156
rect 4187 20154 4243 20156
rect 4267 20154 4323 20156
rect 4347 20154 4403 20156
rect 4107 20102 4153 20154
rect 4153 20102 4163 20154
rect 4187 20102 4217 20154
rect 4217 20102 4229 20154
rect 4229 20102 4243 20154
rect 4267 20102 4281 20154
rect 4281 20102 4293 20154
rect 4293 20102 4323 20154
rect 4347 20102 4357 20154
rect 4357 20102 4403 20154
rect 4107 20100 4163 20102
rect 4187 20100 4243 20102
rect 4267 20100 4323 20102
rect 4347 20100 4403 20102
rect 4107 19066 4163 19068
rect 4187 19066 4243 19068
rect 4267 19066 4323 19068
rect 4347 19066 4403 19068
rect 4107 19014 4153 19066
rect 4153 19014 4163 19066
rect 4187 19014 4217 19066
rect 4217 19014 4229 19066
rect 4229 19014 4243 19066
rect 4267 19014 4281 19066
rect 4281 19014 4293 19066
rect 4293 19014 4323 19066
rect 4347 19014 4357 19066
rect 4357 19014 4403 19066
rect 4107 19012 4163 19014
rect 4187 19012 4243 19014
rect 4267 19012 4323 19014
rect 4347 19012 4403 19014
rect 4767 19610 4823 19612
rect 4847 19610 4903 19612
rect 4927 19610 4983 19612
rect 5007 19610 5063 19612
rect 4767 19558 4813 19610
rect 4813 19558 4823 19610
rect 4847 19558 4877 19610
rect 4877 19558 4889 19610
rect 4889 19558 4903 19610
rect 4927 19558 4941 19610
rect 4941 19558 4953 19610
rect 4953 19558 4983 19610
rect 5007 19558 5017 19610
rect 5017 19558 5063 19610
rect 4767 19556 4823 19558
rect 4847 19556 4903 19558
rect 4927 19556 4983 19558
rect 5007 19556 5063 19558
rect 4802 19352 4858 19408
rect 4767 18522 4823 18524
rect 4847 18522 4903 18524
rect 4927 18522 4983 18524
rect 5007 18522 5063 18524
rect 4767 18470 4813 18522
rect 4813 18470 4823 18522
rect 4847 18470 4877 18522
rect 4877 18470 4889 18522
rect 4889 18470 4903 18522
rect 4927 18470 4941 18522
rect 4941 18470 4953 18522
rect 4953 18470 4983 18522
rect 5007 18470 5017 18522
rect 5017 18470 5063 18522
rect 4767 18468 4823 18470
rect 4847 18468 4903 18470
rect 4927 18468 4983 18470
rect 5007 18468 5063 18470
rect 4107 17978 4163 17980
rect 4187 17978 4243 17980
rect 4267 17978 4323 17980
rect 4347 17978 4403 17980
rect 4107 17926 4153 17978
rect 4153 17926 4163 17978
rect 4187 17926 4217 17978
rect 4217 17926 4229 17978
rect 4229 17926 4243 17978
rect 4267 17926 4281 17978
rect 4281 17926 4293 17978
rect 4293 17926 4323 17978
rect 4347 17926 4357 17978
rect 4357 17926 4403 17978
rect 4107 17924 4163 17926
rect 4187 17924 4243 17926
rect 4267 17924 4323 17926
rect 4347 17924 4403 17926
rect 4107 16890 4163 16892
rect 4187 16890 4243 16892
rect 4267 16890 4323 16892
rect 4347 16890 4403 16892
rect 4107 16838 4153 16890
rect 4153 16838 4163 16890
rect 4187 16838 4217 16890
rect 4217 16838 4229 16890
rect 4229 16838 4243 16890
rect 4267 16838 4281 16890
rect 4281 16838 4293 16890
rect 4293 16838 4323 16890
rect 4347 16838 4357 16890
rect 4357 16838 4403 16890
rect 4107 16836 4163 16838
rect 4187 16836 4243 16838
rect 4267 16836 4323 16838
rect 4347 16836 4403 16838
rect 4107 15802 4163 15804
rect 4187 15802 4243 15804
rect 4267 15802 4323 15804
rect 4347 15802 4403 15804
rect 4107 15750 4153 15802
rect 4153 15750 4163 15802
rect 4187 15750 4217 15802
rect 4217 15750 4229 15802
rect 4229 15750 4243 15802
rect 4267 15750 4281 15802
rect 4281 15750 4293 15802
rect 4293 15750 4323 15802
rect 4347 15750 4357 15802
rect 4357 15750 4403 15802
rect 4107 15748 4163 15750
rect 4187 15748 4243 15750
rect 4267 15748 4323 15750
rect 4347 15748 4403 15750
rect 4767 17434 4823 17436
rect 4847 17434 4903 17436
rect 4927 17434 4983 17436
rect 5007 17434 5063 17436
rect 4767 17382 4813 17434
rect 4813 17382 4823 17434
rect 4847 17382 4877 17434
rect 4877 17382 4889 17434
rect 4889 17382 4903 17434
rect 4927 17382 4941 17434
rect 4941 17382 4953 17434
rect 4953 17382 4983 17434
rect 5007 17382 5017 17434
rect 5017 17382 5063 17434
rect 4767 17380 4823 17382
rect 4847 17380 4903 17382
rect 4927 17380 4983 17382
rect 5007 17380 5063 17382
rect 4767 16346 4823 16348
rect 4847 16346 4903 16348
rect 4927 16346 4983 16348
rect 5007 16346 5063 16348
rect 4767 16294 4813 16346
rect 4813 16294 4823 16346
rect 4847 16294 4877 16346
rect 4877 16294 4889 16346
rect 4889 16294 4903 16346
rect 4927 16294 4941 16346
rect 4941 16294 4953 16346
rect 4953 16294 4983 16346
rect 5007 16294 5017 16346
rect 5017 16294 5063 16346
rect 4767 16292 4823 16294
rect 4847 16292 4903 16294
rect 4927 16292 4983 16294
rect 5007 16292 5063 16294
rect 4767 15258 4823 15260
rect 4847 15258 4903 15260
rect 4927 15258 4983 15260
rect 5007 15258 5063 15260
rect 4767 15206 4813 15258
rect 4813 15206 4823 15258
rect 4847 15206 4877 15258
rect 4877 15206 4889 15258
rect 4889 15206 4903 15258
rect 4927 15206 4941 15258
rect 4941 15206 4953 15258
rect 4953 15206 4983 15258
rect 5007 15206 5017 15258
rect 5017 15206 5063 15258
rect 4767 15204 4823 15206
rect 4847 15204 4903 15206
rect 4927 15204 4983 15206
rect 5007 15204 5063 15206
rect 4107 14714 4163 14716
rect 4187 14714 4243 14716
rect 4267 14714 4323 14716
rect 4347 14714 4403 14716
rect 4107 14662 4153 14714
rect 4153 14662 4163 14714
rect 4187 14662 4217 14714
rect 4217 14662 4229 14714
rect 4229 14662 4243 14714
rect 4267 14662 4281 14714
rect 4281 14662 4293 14714
rect 4293 14662 4323 14714
rect 4347 14662 4357 14714
rect 4357 14662 4403 14714
rect 4107 14660 4163 14662
rect 4187 14660 4243 14662
rect 4267 14660 4323 14662
rect 4347 14660 4403 14662
rect 4107 13626 4163 13628
rect 4187 13626 4243 13628
rect 4267 13626 4323 13628
rect 4347 13626 4403 13628
rect 4107 13574 4153 13626
rect 4153 13574 4163 13626
rect 4187 13574 4217 13626
rect 4217 13574 4229 13626
rect 4229 13574 4243 13626
rect 4267 13574 4281 13626
rect 4281 13574 4293 13626
rect 4293 13574 4323 13626
rect 4347 13574 4357 13626
rect 4357 13574 4403 13626
rect 4107 13572 4163 13574
rect 4187 13572 4243 13574
rect 4267 13572 4323 13574
rect 4347 13572 4403 13574
rect 4107 12538 4163 12540
rect 4187 12538 4243 12540
rect 4267 12538 4323 12540
rect 4347 12538 4403 12540
rect 4107 12486 4153 12538
rect 4153 12486 4163 12538
rect 4187 12486 4217 12538
rect 4217 12486 4229 12538
rect 4229 12486 4243 12538
rect 4267 12486 4281 12538
rect 4281 12486 4293 12538
rect 4293 12486 4323 12538
rect 4347 12486 4357 12538
rect 4357 12486 4403 12538
rect 4107 12484 4163 12486
rect 4187 12484 4243 12486
rect 4267 12484 4323 12486
rect 4347 12484 4403 12486
rect 4342 12164 4398 12200
rect 4342 12144 4344 12164
rect 4344 12144 4396 12164
rect 4396 12144 4398 12164
rect 4107 11450 4163 11452
rect 4187 11450 4243 11452
rect 4267 11450 4323 11452
rect 4347 11450 4403 11452
rect 4107 11398 4153 11450
rect 4153 11398 4163 11450
rect 4187 11398 4217 11450
rect 4217 11398 4229 11450
rect 4229 11398 4243 11450
rect 4267 11398 4281 11450
rect 4281 11398 4293 11450
rect 4293 11398 4323 11450
rect 4347 11398 4357 11450
rect 4357 11398 4403 11450
rect 4107 11396 4163 11398
rect 4187 11396 4243 11398
rect 4267 11396 4323 11398
rect 4347 11396 4403 11398
rect 4107 10362 4163 10364
rect 4187 10362 4243 10364
rect 4267 10362 4323 10364
rect 4347 10362 4403 10364
rect 4107 10310 4153 10362
rect 4153 10310 4163 10362
rect 4187 10310 4217 10362
rect 4217 10310 4229 10362
rect 4229 10310 4243 10362
rect 4267 10310 4281 10362
rect 4281 10310 4293 10362
rect 4293 10310 4323 10362
rect 4347 10310 4357 10362
rect 4357 10310 4403 10362
rect 4107 10308 4163 10310
rect 4187 10308 4243 10310
rect 4267 10308 4323 10310
rect 4347 10308 4403 10310
rect 4767 14170 4823 14172
rect 4847 14170 4903 14172
rect 4927 14170 4983 14172
rect 5007 14170 5063 14172
rect 4767 14118 4813 14170
rect 4813 14118 4823 14170
rect 4847 14118 4877 14170
rect 4877 14118 4889 14170
rect 4889 14118 4903 14170
rect 4927 14118 4941 14170
rect 4941 14118 4953 14170
rect 4953 14118 4983 14170
rect 5007 14118 5017 14170
rect 5017 14118 5063 14170
rect 4767 14116 4823 14118
rect 4847 14116 4903 14118
rect 4927 14116 4983 14118
rect 5007 14116 5063 14118
rect 4767 13082 4823 13084
rect 4847 13082 4903 13084
rect 4927 13082 4983 13084
rect 5007 13082 5063 13084
rect 4767 13030 4813 13082
rect 4813 13030 4823 13082
rect 4847 13030 4877 13082
rect 4877 13030 4889 13082
rect 4889 13030 4903 13082
rect 4927 13030 4941 13082
rect 4941 13030 4953 13082
rect 4953 13030 4983 13082
rect 5007 13030 5017 13082
rect 5017 13030 5063 13082
rect 4767 13028 4823 13030
rect 4847 13028 4903 13030
rect 4927 13028 4983 13030
rect 5007 13028 5063 13030
rect 4767 11994 4823 11996
rect 4847 11994 4903 11996
rect 4927 11994 4983 11996
rect 5007 11994 5063 11996
rect 4767 11942 4813 11994
rect 4813 11942 4823 11994
rect 4847 11942 4877 11994
rect 4877 11942 4889 11994
rect 4889 11942 4903 11994
rect 4927 11942 4941 11994
rect 4941 11942 4953 11994
rect 4953 11942 4983 11994
rect 5007 11942 5017 11994
rect 5017 11942 5063 11994
rect 4767 11940 4823 11942
rect 4847 11940 4903 11942
rect 4927 11940 4983 11942
rect 5007 11940 5063 11942
rect 4710 11756 4766 11792
rect 4710 11736 4712 11756
rect 4712 11736 4764 11756
rect 4764 11736 4766 11756
rect 5446 12280 5502 12336
rect 6642 17484 6644 17504
rect 6644 17484 6696 17504
rect 6696 17484 6698 17504
rect 6642 17448 6698 17484
rect 10409 22330 10465 22332
rect 10489 22330 10545 22332
rect 10569 22330 10625 22332
rect 10649 22330 10705 22332
rect 10409 22278 10455 22330
rect 10455 22278 10465 22330
rect 10489 22278 10519 22330
rect 10519 22278 10531 22330
rect 10531 22278 10545 22330
rect 10569 22278 10583 22330
rect 10583 22278 10595 22330
rect 10595 22278 10625 22330
rect 10649 22278 10659 22330
rect 10659 22278 10705 22330
rect 10409 22276 10465 22278
rect 10489 22276 10545 22278
rect 10569 22276 10625 22278
rect 10649 22276 10705 22278
rect 10409 21242 10465 21244
rect 10489 21242 10545 21244
rect 10569 21242 10625 21244
rect 10649 21242 10705 21244
rect 10409 21190 10455 21242
rect 10455 21190 10465 21242
rect 10489 21190 10519 21242
rect 10519 21190 10531 21242
rect 10531 21190 10545 21242
rect 10569 21190 10583 21242
rect 10583 21190 10595 21242
rect 10595 21190 10625 21242
rect 10649 21190 10659 21242
rect 10659 21190 10705 21242
rect 10409 21188 10465 21190
rect 10489 21188 10545 21190
rect 10569 21188 10625 21190
rect 10649 21188 10705 21190
rect 11069 21786 11125 21788
rect 11149 21786 11205 21788
rect 11229 21786 11285 21788
rect 11309 21786 11365 21788
rect 11069 21734 11115 21786
rect 11115 21734 11125 21786
rect 11149 21734 11179 21786
rect 11179 21734 11191 21786
rect 11191 21734 11205 21786
rect 11229 21734 11243 21786
rect 11243 21734 11255 21786
rect 11255 21734 11285 21786
rect 11309 21734 11319 21786
rect 11319 21734 11365 21786
rect 11069 21732 11125 21734
rect 11149 21732 11205 21734
rect 11229 21732 11285 21734
rect 11309 21732 11365 21734
rect 7930 17856 7986 17912
rect 5630 12280 5686 12336
rect 5354 11736 5410 11792
rect 5538 11772 5540 11792
rect 5540 11772 5592 11792
rect 5592 11772 5594 11792
rect 5538 11736 5594 11772
rect 5630 11600 5686 11656
rect 5538 11228 5540 11248
rect 5540 11228 5592 11248
rect 5592 11228 5594 11248
rect 5538 11192 5594 11228
rect 6366 11228 6368 11248
rect 6368 11228 6420 11248
rect 6420 11228 6422 11248
rect 6366 11192 6422 11228
rect 6274 11056 6330 11112
rect 6826 12144 6882 12200
rect 6734 11756 6790 11792
rect 6734 11736 6736 11756
rect 6736 11736 6788 11756
rect 6788 11736 6790 11756
rect 6734 11600 6790 11656
rect 4767 10906 4823 10908
rect 4847 10906 4903 10908
rect 4927 10906 4983 10908
rect 5007 10906 5063 10908
rect 4767 10854 4813 10906
rect 4813 10854 4823 10906
rect 4847 10854 4877 10906
rect 4877 10854 4889 10906
rect 4889 10854 4903 10906
rect 4927 10854 4941 10906
rect 4941 10854 4953 10906
rect 4953 10854 4983 10906
rect 5007 10854 5017 10906
rect 5017 10854 5063 10906
rect 4767 10852 4823 10854
rect 4847 10852 4903 10854
rect 4927 10852 4983 10854
rect 5007 10852 5063 10854
rect 4767 9818 4823 9820
rect 4847 9818 4903 9820
rect 4927 9818 4983 9820
rect 5007 9818 5063 9820
rect 4767 9766 4813 9818
rect 4813 9766 4823 9818
rect 4847 9766 4877 9818
rect 4877 9766 4889 9818
rect 4889 9766 4903 9818
rect 4927 9766 4941 9818
rect 4941 9766 4953 9818
rect 4953 9766 4983 9818
rect 5007 9766 5017 9818
rect 5017 9766 5063 9818
rect 4767 9764 4823 9766
rect 4847 9764 4903 9766
rect 4927 9764 4983 9766
rect 5007 9764 5063 9766
rect 4107 9274 4163 9276
rect 4187 9274 4243 9276
rect 4267 9274 4323 9276
rect 4347 9274 4403 9276
rect 4107 9222 4153 9274
rect 4153 9222 4163 9274
rect 4187 9222 4217 9274
rect 4217 9222 4229 9274
rect 4229 9222 4243 9274
rect 4267 9222 4281 9274
rect 4281 9222 4293 9274
rect 4293 9222 4323 9274
rect 4347 9222 4357 9274
rect 4357 9222 4403 9274
rect 4107 9220 4163 9222
rect 4187 9220 4243 9222
rect 4267 9220 4323 9222
rect 4347 9220 4403 9222
rect 4802 9052 4804 9072
rect 4804 9052 4856 9072
rect 4856 9052 4858 9072
rect 4802 9016 4858 9052
rect 4894 8880 4950 8936
rect 4767 8730 4823 8732
rect 4847 8730 4903 8732
rect 4927 8730 4983 8732
rect 5007 8730 5063 8732
rect 4767 8678 4813 8730
rect 4813 8678 4823 8730
rect 4847 8678 4877 8730
rect 4877 8678 4889 8730
rect 4889 8678 4903 8730
rect 4927 8678 4941 8730
rect 4941 8678 4953 8730
rect 4953 8678 4983 8730
rect 5007 8678 5017 8730
rect 5017 8678 5063 8730
rect 4767 8676 4823 8678
rect 4847 8676 4903 8678
rect 4927 8676 4983 8678
rect 5007 8676 5063 8678
rect 4107 8186 4163 8188
rect 4187 8186 4243 8188
rect 4267 8186 4323 8188
rect 4347 8186 4403 8188
rect 4107 8134 4153 8186
rect 4153 8134 4163 8186
rect 4187 8134 4217 8186
rect 4217 8134 4229 8186
rect 4229 8134 4243 8186
rect 4267 8134 4281 8186
rect 4281 8134 4293 8186
rect 4293 8134 4323 8186
rect 4347 8134 4357 8186
rect 4357 8134 4403 8186
rect 4107 8132 4163 8134
rect 4187 8132 4243 8134
rect 4267 8132 4323 8134
rect 4347 8132 4403 8134
rect 4986 8472 5042 8528
rect 4767 7642 4823 7644
rect 4847 7642 4903 7644
rect 4927 7642 4983 7644
rect 5007 7642 5063 7644
rect 4767 7590 4813 7642
rect 4813 7590 4823 7642
rect 4847 7590 4877 7642
rect 4877 7590 4889 7642
rect 4889 7590 4903 7642
rect 4927 7590 4941 7642
rect 4941 7590 4953 7642
rect 4953 7590 4983 7642
rect 5007 7590 5017 7642
rect 5017 7590 5063 7642
rect 4767 7588 4823 7590
rect 4847 7588 4903 7590
rect 4927 7588 4983 7590
rect 5007 7588 5063 7590
rect 4107 7098 4163 7100
rect 4187 7098 4243 7100
rect 4267 7098 4323 7100
rect 4347 7098 4403 7100
rect 4107 7046 4153 7098
rect 4153 7046 4163 7098
rect 4187 7046 4217 7098
rect 4217 7046 4229 7098
rect 4229 7046 4243 7098
rect 4267 7046 4281 7098
rect 4281 7046 4293 7098
rect 4293 7046 4323 7098
rect 4347 7046 4357 7098
rect 4357 7046 4403 7098
rect 4107 7044 4163 7046
rect 4187 7044 4243 7046
rect 4267 7044 4323 7046
rect 4347 7044 4403 7046
rect 4767 6554 4823 6556
rect 4847 6554 4903 6556
rect 4927 6554 4983 6556
rect 5007 6554 5063 6556
rect 4767 6502 4813 6554
rect 4813 6502 4823 6554
rect 4847 6502 4877 6554
rect 4877 6502 4889 6554
rect 4889 6502 4903 6554
rect 4927 6502 4941 6554
rect 4941 6502 4953 6554
rect 4953 6502 4983 6554
rect 5007 6502 5017 6554
rect 5017 6502 5063 6554
rect 4767 6500 4823 6502
rect 4847 6500 4903 6502
rect 4927 6500 4983 6502
rect 5007 6500 5063 6502
rect 4107 6010 4163 6012
rect 4187 6010 4243 6012
rect 4267 6010 4323 6012
rect 4347 6010 4403 6012
rect 4107 5958 4153 6010
rect 4153 5958 4163 6010
rect 4187 5958 4217 6010
rect 4217 5958 4229 6010
rect 4229 5958 4243 6010
rect 4267 5958 4281 6010
rect 4281 5958 4293 6010
rect 4293 5958 4323 6010
rect 4347 5958 4357 6010
rect 4357 5958 4403 6010
rect 4107 5956 4163 5958
rect 4187 5956 4243 5958
rect 4267 5956 4323 5958
rect 4347 5956 4403 5958
rect 5538 8608 5594 8664
rect 5630 8064 5686 8120
rect 4767 5466 4823 5468
rect 4847 5466 4903 5468
rect 4927 5466 4983 5468
rect 5007 5466 5063 5468
rect 4767 5414 4813 5466
rect 4813 5414 4823 5466
rect 4847 5414 4877 5466
rect 4877 5414 4889 5466
rect 4889 5414 4903 5466
rect 4927 5414 4941 5466
rect 4941 5414 4953 5466
rect 4953 5414 4983 5466
rect 5007 5414 5017 5466
rect 5017 5414 5063 5466
rect 4767 5412 4823 5414
rect 4847 5412 4903 5414
rect 4927 5412 4983 5414
rect 5007 5412 5063 5414
rect 4107 4922 4163 4924
rect 4187 4922 4243 4924
rect 4267 4922 4323 4924
rect 4347 4922 4403 4924
rect 4107 4870 4153 4922
rect 4153 4870 4163 4922
rect 4187 4870 4217 4922
rect 4217 4870 4229 4922
rect 4229 4870 4243 4922
rect 4267 4870 4281 4922
rect 4281 4870 4293 4922
rect 4293 4870 4323 4922
rect 4347 4870 4357 4922
rect 4357 4870 4403 4922
rect 4107 4868 4163 4870
rect 4187 4868 4243 4870
rect 4267 4868 4323 4870
rect 4347 4868 4403 4870
rect 6458 9036 6514 9072
rect 6458 9016 6460 9036
rect 6460 9016 6512 9036
rect 6512 9016 6514 9036
rect 11069 20698 11125 20700
rect 11149 20698 11205 20700
rect 11229 20698 11285 20700
rect 11309 20698 11365 20700
rect 11069 20646 11115 20698
rect 11115 20646 11125 20698
rect 11149 20646 11179 20698
rect 11179 20646 11191 20698
rect 11191 20646 11205 20698
rect 11229 20646 11243 20698
rect 11243 20646 11255 20698
rect 11255 20646 11285 20698
rect 11309 20646 11319 20698
rect 11319 20646 11365 20698
rect 11069 20644 11125 20646
rect 11149 20644 11205 20646
rect 11229 20644 11285 20646
rect 11309 20644 11365 20646
rect 10409 20154 10465 20156
rect 10489 20154 10545 20156
rect 10569 20154 10625 20156
rect 10649 20154 10705 20156
rect 10409 20102 10455 20154
rect 10455 20102 10465 20154
rect 10489 20102 10519 20154
rect 10519 20102 10531 20154
rect 10531 20102 10545 20154
rect 10569 20102 10583 20154
rect 10583 20102 10595 20154
rect 10595 20102 10625 20154
rect 10649 20102 10659 20154
rect 10659 20102 10705 20154
rect 10409 20100 10465 20102
rect 10489 20100 10545 20102
rect 10569 20100 10625 20102
rect 10649 20100 10705 20102
rect 11069 19610 11125 19612
rect 11149 19610 11205 19612
rect 11229 19610 11285 19612
rect 11309 19610 11365 19612
rect 11069 19558 11115 19610
rect 11115 19558 11125 19610
rect 11149 19558 11179 19610
rect 11179 19558 11191 19610
rect 11191 19558 11205 19610
rect 11229 19558 11243 19610
rect 11243 19558 11255 19610
rect 11255 19558 11285 19610
rect 11309 19558 11319 19610
rect 11319 19558 11365 19610
rect 11069 19556 11125 19558
rect 11149 19556 11205 19558
rect 11229 19556 11285 19558
rect 11309 19556 11365 19558
rect 10322 19352 10378 19408
rect 10409 19066 10465 19068
rect 10489 19066 10545 19068
rect 10569 19066 10625 19068
rect 10649 19066 10705 19068
rect 10409 19014 10455 19066
rect 10455 19014 10465 19066
rect 10489 19014 10519 19066
rect 10519 19014 10531 19066
rect 10531 19014 10545 19066
rect 10569 19014 10583 19066
rect 10583 19014 10595 19066
rect 10595 19014 10625 19066
rect 10649 19014 10659 19066
rect 10659 19014 10705 19066
rect 10409 19012 10465 19014
rect 10489 19012 10545 19014
rect 10569 19012 10625 19014
rect 10649 19012 10705 19014
rect 11069 18522 11125 18524
rect 11149 18522 11205 18524
rect 11229 18522 11285 18524
rect 11309 18522 11365 18524
rect 11069 18470 11115 18522
rect 11115 18470 11125 18522
rect 11149 18470 11179 18522
rect 11179 18470 11191 18522
rect 11191 18470 11205 18522
rect 11229 18470 11243 18522
rect 11243 18470 11255 18522
rect 11255 18470 11285 18522
rect 11309 18470 11319 18522
rect 11319 18470 11365 18522
rect 11069 18468 11125 18470
rect 11149 18468 11205 18470
rect 11229 18468 11285 18470
rect 11309 18468 11365 18470
rect 10138 17856 10194 17912
rect 10409 17978 10465 17980
rect 10489 17978 10545 17980
rect 10569 17978 10625 17980
rect 10649 17978 10705 17980
rect 10409 17926 10455 17978
rect 10455 17926 10465 17978
rect 10489 17926 10519 17978
rect 10519 17926 10531 17978
rect 10531 17926 10545 17978
rect 10569 17926 10583 17978
rect 10583 17926 10595 17978
rect 10595 17926 10625 17978
rect 10649 17926 10659 17978
rect 10659 17926 10705 17978
rect 10409 17924 10465 17926
rect 10489 17924 10545 17926
rect 10569 17924 10625 17926
rect 10649 17924 10705 17926
rect 10409 16890 10465 16892
rect 10489 16890 10545 16892
rect 10569 16890 10625 16892
rect 10649 16890 10705 16892
rect 10409 16838 10455 16890
rect 10455 16838 10465 16890
rect 10489 16838 10519 16890
rect 10519 16838 10531 16890
rect 10531 16838 10545 16890
rect 10569 16838 10583 16890
rect 10583 16838 10595 16890
rect 10595 16838 10625 16890
rect 10649 16838 10659 16890
rect 10659 16838 10705 16890
rect 10409 16836 10465 16838
rect 10489 16836 10545 16838
rect 10569 16836 10625 16838
rect 10649 16836 10705 16838
rect 11069 17434 11125 17436
rect 11149 17434 11205 17436
rect 11229 17434 11285 17436
rect 11309 17434 11365 17436
rect 11069 17382 11115 17434
rect 11115 17382 11125 17434
rect 11149 17382 11179 17434
rect 11179 17382 11191 17434
rect 11191 17382 11205 17434
rect 11229 17382 11243 17434
rect 11243 17382 11255 17434
rect 11255 17382 11285 17434
rect 11309 17382 11319 17434
rect 11319 17382 11365 17434
rect 11069 17380 11125 17382
rect 11149 17380 11205 17382
rect 11229 17380 11285 17382
rect 11309 17380 11365 17382
rect 16711 26682 16767 26684
rect 16791 26682 16847 26684
rect 16871 26682 16927 26684
rect 16951 26682 17007 26684
rect 16711 26630 16757 26682
rect 16757 26630 16767 26682
rect 16791 26630 16821 26682
rect 16821 26630 16833 26682
rect 16833 26630 16847 26682
rect 16871 26630 16885 26682
rect 16885 26630 16897 26682
rect 16897 26630 16927 26682
rect 16951 26630 16961 26682
rect 16961 26630 17007 26682
rect 16711 26628 16767 26630
rect 16791 26628 16847 26630
rect 16871 26628 16927 26630
rect 16951 26628 17007 26630
rect 14278 20884 14280 20904
rect 14280 20884 14332 20904
rect 14332 20884 14334 20904
rect 11069 16346 11125 16348
rect 11149 16346 11205 16348
rect 11229 16346 11285 16348
rect 11309 16346 11365 16348
rect 11069 16294 11115 16346
rect 11115 16294 11125 16346
rect 11149 16294 11179 16346
rect 11179 16294 11191 16346
rect 11191 16294 11205 16346
rect 11229 16294 11243 16346
rect 11243 16294 11255 16346
rect 11255 16294 11285 16346
rect 11309 16294 11319 16346
rect 11319 16294 11365 16346
rect 11069 16292 11125 16294
rect 11149 16292 11205 16294
rect 11229 16292 11285 16294
rect 11309 16292 11365 16294
rect 10409 15802 10465 15804
rect 10489 15802 10545 15804
rect 10569 15802 10625 15804
rect 10649 15802 10705 15804
rect 10409 15750 10455 15802
rect 10455 15750 10465 15802
rect 10489 15750 10519 15802
rect 10519 15750 10531 15802
rect 10531 15750 10545 15802
rect 10569 15750 10583 15802
rect 10583 15750 10595 15802
rect 10595 15750 10625 15802
rect 10649 15750 10659 15802
rect 10659 15750 10705 15802
rect 10409 15748 10465 15750
rect 10489 15748 10545 15750
rect 10569 15748 10625 15750
rect 10649 15748 10705 15750
rect 8206 12144 8262 12200
rect 7654 11056 7710 11112
rect 11069 15258 11125 15260
rect 11149 15258 11205 15260
rect 11229 15258 11285 15260
rect 11309 15258 11365 15260
rect 11069 15206 11115 15258
rect 11115 15206 11125 15258
rect 11149 15206 11179 15258
rect 11179 15206 11191 15258
rect 11191 15206 11205 15258
rect 11229 15206 11243 15258
rect 11243 15206 11255 15258
rect 11255 15206 11285 15258
rect 11309 15206 11319 15258
rect 11319 15206 11365 15258
rect 11069 15204 11125 15206
rect 11149 15204 11205 15206
rect 11229 15204 11285 15206
rect 11309 15204 11365 15206
rect 10409 14714 10465 14716
rect 10489 14714 10545 14716
rect 10569 14714 10625 14716
rect 10649 14714 10705 14716
rect 10409 14662 10455 14714
rect 10455 14662 10465 14714
rect 10489 14662 10519 14714
rect 10519 14662 10531 14714
rect 10531 14662 10545 14714
rect 10569 14662 10583 14714
rect 10583 14662 10595 14714
rect 10595 14662 10625 14714
rect 10649 14662 10659 14714
rect 10659 14662 10705 14714
rect 10409 14660 10465 14662
rect 10489 14660 10545 14662
rect 10569 14660 10625 14662
rect 10649 14660 10705 14662
rect 4767 4378 4823 4380
rect 4847 4378 4903 4380
rect 4927 4378 4983 4380
rect 5007 4378 5063 4380
rect 4767 4326 4813 4378
rect 4813 4326 4823 4378
rect 4847 4326 4877 4378
rect 4877 4326 4889 4378
rect 4889 4326 4903 4378
rect 4927 4326 4941 4378
rect 4941 4326 4953 4378
rect 4953 4326 4983 4378
rect 5007 4326 5017 4378
rect 5017 4326 5063 4378
rect 4767 4324 4823 4326
rect 4847 4324 4903 4326
rect 4927 4324 4983 4326
rect 5007 4324 5063 4326
rect 3698 4120 3754 4176
rect 4107 3834 4163 3836
rect 4187 3834 4243 3836
rect 4267 3834 4323 3836
rect 4347 3834 4403 3836
rect 4107 3782 4153 3834
rect 4153 3782 4163 3834
rect 4187 3782 4217 3834
rect 4217 3782 4229 3834
rect 4229 3782 4243 3834
rect 4267 3782 4281 3834
rect 4281 3782 4293 3834
rect 4293 3782 4323 3834
rect 4347 3782 4357 3834
rect 4357 3782 4403 3834
rect 4107 3780 4163 3782
rect 4187 3780 4243 3782
rect 4267 3780 4323 3782
rect 4347 3780 4403 3782
rect 4894 3476 4896 3496
rect 4896 3476 4948 3496
rect 4948 3476 4950 3496
rect 4894 3440 4950 3476
rect 4767 3290 4823 3292
rect 4847 3290 4903 3292
rect 4927 3290 4983 3292
rect 5007 3290 5063 3292
rect 4767 3238 4813 3290
rect 4813 3238 4823 3290
rect 4847 3238 4877 3290
rect 4877 3238 4889 3290
rect 4889 3238 4903 3290
rect 4927 3238 4941 3290
rect 4941 3238 4953 3290
rect 4953 3238 4983 3290
rect 5007 3238 5017 3290
rect 5017 3238 5063 3290
rect 4767 3236 4823 3238
rect 4847 3236 4903 3238
rect 4927 3236 4983 3238
rect 5007 3236 5063 3238
rect 4107 2746 4163 2748
rect 4187 2746 4243 2748
rect 4267 2746 4323 2748
rect 4347 2746 4403 2748
rect 4107 2694 4153 2746
rect 4153 2694 4163 2746
rect 4187 2694 4217 2746
rect 4217 2694 4229 2746
rect 4229 2694 4243 2746
rect 4267 2694 4281 2746
rect 4281 2694 4293 2746
rect 4293 2694 4323 2746
rect 4347 2694 4357 2746
rect 4357 2694 4403 2746
rect 4107 2692 4163 2694
rect 4187 2692 4243 2694
rect 4267 2692 4323 2694
rect 4347 2692 4403 2694
rect 7470 3440 7526 3496
rect 10409 13626 10465 13628
rect 10489 13626 10545 13628
rect 10569 13626 10625 13628
rect 10649 13626 10705 13628
rect 10409 13574 10455 13626
rect 10455 13574 10465 13626
rect 10489 13574 10519 13626
rect 10519 13574 10531 13626
rect 10531 13574 10545 13626
rect 10569 13574 10583 13626
rect 10583 13574 10595 13626
rect 10595 13574 10625 13626
rect 10649 13574 10659 13626
rect 10659 13574 10705 13626
rect 10409 13572 10465 13574
rect 10489 13572 10545 13574
rect 10569 13572 10625 13574
rect 10649 13572 10705 13574
rect 10409 12538 10465 12540
rect 10489 12538 10545 12540
rect 10569 12538 10625 12540
rect 10649 12538 10705 12540
rect 10409 12486 10455 12538
rect 10455 12486 10465 12538
rect 10489 12486 10519 12538
rect 10519 12486 10531 12538
rect 10531 12486 10545 12538
rect 10569 12486 10583 12538
rect 10583 12486 10595 12538
rect 10595 12486 10625 12538
rect 10649 12486 10659 12538
rect 10659 12486 10705 12538
rect 10409 12484 10465 12486
rect 10489 12484 10545 12486
rect 10569 12484 10625 12486
rect 10649 12484 10705 12486
rect 11069 14170 11125 14172
rect 11149 14170 11205 14172
rect 11229 14170 11285 14172
rect 11309 14170 11365 14172
rect 11069 14118 11115 14170
rect 11115 14118 11125 14170
rect 11149 14118 11179 14170
rect 11179 14118 11191 14170
rect 11191 14118 11205 14170
rect 11229 14118 11243 14170
rect 11243 14118 11255 14170
rect 11255 14118 11285 14170
rect 11309 14118 11319 14170
rect 11319 14118 11365 14170
rect 11069 14116 11125 14118
rect 11149 14116 11205 14118
rect 11229 14116 11285 14118
rect 11309 14116 11365 14118
rect 11069 13082 11125 13084
rect 11149 13082 11205 13084
rect 11229 13082 11285 13084
rect 11309 13082 11365 13084
rect 11069 13030 11115 13082
rect 11115 13030 11125 13082
rect 11149 13030 11179 13082
rect 11179 13030 11191 13082
rect 11191 13030 11205 13082
rect 11229 13030 11243 13082
rect 11243 13030 11255 13082
rect 11255 13030 11285 13082
rect 11309 13030 11319 13082
rect 11319 13030 11365 13082
rect 11069 13028 11125 13030
rect 11149 13028 11205 13030
rect 11229 13028 11285 13030
rect 11309 13028 11365 13030
rect 10409 11450 10465 11452
rect 10489 11450 10545 11452
rect 10569 11450 10625 11452
rect 10649 11450 10705 11452
rect 10409 11398 10455 11450
rect 10455 11398 10465 11450
rect 10489 11398 10519 11450
rect 10519 11398 10531 11450
rect 10531 11398 10545 11450
rect 10569 11398 10583 11450
rect 10583 11398 10595 11450
rect 10595 11398 10625 11450
rect 10649 11398 10659 11450
rect 10659 11398 10705 11450
rect 10409 11396 10465 11398
rect 10489 11396 10545 11398
rect 10569 11396 10625 11398
rect 10649 11396 10705 11398
rect 11069 11994 11125 11996
rect 11149 11994 11205 11996
rect 11229 11994 11285 11996
rect 11309 11994 11365 11996
rect 11069 11942 11115 11994
rect 11115 11942 11125 11994
rect 11149 11942 11179 11994
rect 11179 11942 11191 11994
rect 11191 11942 11205 11994
rect 11229 11942 11243 11994
rect 11243 11942 11255 11994
rect 11255 11942 11285 11994
rect 11309 11942 11319 11994
rect 11319 11942 11365 11994
rect 11069 11940 11125 11942
rect 11149 11940 11205 11942
rect 11229 11940 11285 11942
rect 11309 11940 11365 11942
rect 10409 10362 10465 10364
rect 10489 10362 10545 10364
rect 10569 10362 10625 10364
rect 10649 10362 10705 10364
rect 10409 10310 10455 10362
rect 10455 10310 10465 10362
rect 10489 10310 10519 10362
rect 10519 10310 10531 10362
rect 10531 10310 10545 10362
rect 10569 10310 10583 10362
rect 10583 10310 10595 10362
rect 10595 10310 10625 10362
rect 10649 10310 10659 10362
rect 10659 10310 10705 10362
rect 10409 10308 10465 10310
rect 10489 10308 10545 10310
rect 10569 10308 10625 10310
rect 10649 10308 10705 10310
rect 11069 10906 11125 10908
rect 11149 10906 11205 10908
rect 11229 10906 11285 10908
rect 11309 10906 11365 10908
rect 11069 10854 11115 10906
rect 11115 10854 11125 10906
rect 11149 10854 11179 10906
rect 11179 10854 11191 10906
rect 11191 10854 11205 10906
rect 11229 10854 11243 10906
rect 11243 10854 11255 10906
rect 11255 10854 11285 10906
rect 11309 10854 11319 10906
rect 11319 10854 11365 10906
rect 11069 10852 11125 10854
rect 11149 10852 11205 10854
rect 11229 10852 11285 10854
rect 11309 10852 11365 10854
rect 10409 9274 10465 9276
rect 10489 9274 10545 9276
rect 10569 9274 10625 9276
rect 10649 9274 10705 9276
rect 10409 9222 10455 9274
rect 10455 9222 10465 9274
rect 10489 9222 10519 9274
rect 10519 9222 10531 9274
rect 10531 9222 10545 9274
rect 10569 9222 10583 9274
rect 10583 9222 10595 9274
rect 10595 9222 10625 9274
rect 10649 9222 10659 9274
rect 10659 9222 10705 9274
rect 10409 9220 10465 9222
rect 10489 9220 10545 9222
rect 10569 9220 10625 9222
rect 10649 9220 10705 9222
rect 11069 9818 11125 9820
rect 11149 9818 11205 9820
rect 11229 9818 11285 9820
rect 11309 9818 11365 9820
rect 11069 9766 11115 9818
rect 11115 9766 11125 9818
rect 11149 9766 11179 9818
rect 11179 9766 11191 9818
rect 11191 9766 11205 9818
rect 11229 9766 11243 9818
rect 11243 9766 11255 9818
rect 11255 9766 11285 9818
rect 11309 9766 11319 9818
rect 11319 9766 11365 9818
rect 11069 9764 11125 9766
rect 11149 9764 11205 9766
rect 11229 9764 11285 9766
rect 11309 9764 11365 9766
rect 11069 8730 11125 8732
rect 11149 8730 11205 8732
rect 11229 8730 11285 8732
rect 11309 8730 11365 8732
rect 11069 8678 11115 8730
rect 11115 8678 11125 8730
rect 11149 8678 11179 8730
rect 11179 8678 11191 8730
rect 11191 8678 11205 8730
rect 11229 8678 11243 8730
rect 11243 8678 11255 8730
rect 11255 8678 11285 8730
rect 11309 8678 11319 8730
rect 11319 8678 11365 8730
rect 11069 8676 11125 8678
rect 11149 8676 11205 8678
rect 11229 8676 11285 8678
rect 11309 8676 11365 8678
rect 10409 8186 10465 8188
rect 10489 8186 10545 8188
rect 10569 8186 10625 8188
rect 10649 8186 10705 8188
rect 10409 8134 10455 8186
rect 10455 8134 10465 8186
rect 10489 8134 10519 8186
rect 10519 8134 10531 8186
rect 10531 8134 10545 8186
rect 10569 8134 10583 8186
rect 10583 8134 10595 8186
rect 10595 8134 10625 8186
rect 10649 8134 10659 8186
rect 10659 8134 10705 8186
rect 10409 8132 10465 8134
rect 10489 8132 10545 8134
rect 10569 8132 10625 8134
rect 10649 8132 10705 8134
rect 10409 7098 10465 7100
rect 10489 7098 10545 7100
rect 10569 7098 10625 7100
rect 10649 7098 10705 7100
rect 10409 7046 10455 7098
rect 10455 7046 10465 7098
rect 10489 7046 10519 7098
rect 10519 7046 10531 7098
rect 10531 7046 10545 7098
rect 10569 7046 10583 7098
rect 10583 7046 10595 7098
rect 10595 7046 10625 7098
rect 10649 7046 10659 7098
rect 10659 7046 10705 7098
rect 10409 7044 10465 7046
rect 10489 7044 10545 7046
rect 10569 7044 10625 7046
rect 10649 7044 10705 7046
rect 10409 6010 10465 6012
rect 10489 6010 10545 6012
rect 10569 6010 10625 6012
rect 10649 6010 10705 6012
rect 10409 5958 10455 6010
rect 10455 5958 10465 6010
rect 10489 5958 10519 6010
rect 10519 5958 10531 6010
rect 10531 5958 10545 6010
rect 10569 5958 10583 6010
rect 10583 5958 10595 6010
rect 10595 5958 10625 6010
rect 10649 5958 10659 6010
rect 10659 5958 10705 6010
rect 10409 5956 10465 5958
rect 10489 5956 10545 5958
rect 10569 5956 10625 5958
rect 10649 5956 10705 5958
rect 10409 4922 10465 4924
rect 10489 4922 10545 4924
rect 10569 4922 10625 4924
rect 10649 4922 10705 4924
rect 10409 4870 10455 4922
rect 10455 4870 10465 4922
rect 10489 4870 10519 4922
rect 10519 4870 10531 4922
rect 10531 4870 10545 4922
rect 10569 4870 10583 4922
rect 10583 4870 10595 4922
rect 10595 4870 10625 4922
rect 10649 4870 10659 4922
rect 10659 4870 10705 4922
rect 10409 4868 10465 4870
rect 10489 4868 10545 4870
rect 10569 4868 10625 4870
rect 10649 4868 10705 4870
rect 10409 3834 10465 3836
rect 10489 3834 10545 3836
rect 10569 3834 10625 3836
rect 10649 3834 10705 3836
rect 10409 3782 10455 3834
rect 10455 3782 10465 3834
rect 10489 3782 10519 3834
rect 10519 3782 10531 3834
rect 10531 3782 10545 3834
rect 10569 3782 10583 3834
rect 10583 3782 10595 3834
rect 10595 3782 10625 3834
rect 10649 3782 10659 3834
rect 10659 3782 10705 3834
rect 10409 3780 10465 3782
rect 10489 3780 10545 3782
rect 10569 3780 10625 3782
rect 10649 3780 10705 3782
rect 10409 2746 10465 2748
rect 10489 2746 10545 2748
rect 10569 2746 10625 2748
rect 10649 2746 10705 2748
rect 10409 2694 10455 2746
rect 10455 2694 10465 2746
rect 10489 2694 10519 2746
rect 10519 2694 10531 2746
rect 10531 2694 10545 2746
rect 10569 2694 10583 2746
rect 10583 2694 10595 2746
rect 10595 2694 10625 2746
rect 10649 2694 10659 2746
rect 10659 2694 10705 2746
rect 10409 2692 10465 2694
rect 10489 2692 10545 2694
rect 10569 2692 10625 2694
rect 10649 2692 10705 2694
rect 4767 2202 4823 2204
rect 4847 2202 4903 2204
rect 4927 2202 4983 2204
rect 5007 2202 5063 2204
rect 4767 2150 4813 2202
rect 4813 2150 4823 2202
rect 4847 2150 4877 2202
rect 4877 2150 4889 2202
rect 4889 2150 4903 2202
rect 4927 2150 4941 2202
rect 4941 2150 4953 2202
rect 4953 2150 4983 2202
rect 5007 2150 5017 2202
rect 5017 2150 5063 2202
rect 4767 2148 4823 2150
rect 4847 2148 4903 2150
rect 4927 2148 4983 2150
rect 5007 2148 5063 2150
rect 11069 7642 11125 7644
rect 11149 7642 11205 7644
rect 11229 7642 11285 7644
rect 11309 7642 11365 7644
rect 11069 7590 11115 7642
rect 11115 7590 11125 7642
rect 11149 7590 11179 7642
rect 11179 7590 11191 7642
rect 11191 7590 11205 7642
rect 11229 7590 11243 7642
rect 11243 7590 11255 7642
rect 11255 7590 11285 7642
rect 11309 7590 11319 7642
rect 11319 7590 11365 7642
rect 11069 7588 11125 7590
rect 11149 7588 11205 7590
rect 11229 7588 11285 7590
rect 11309 7588 11365 7590
rect 11069 6554 11125 6556
rect 11149 6554 11205 6556
rect 11229 6554 11285 6556
rect 11309 6554 11365 6556
rect 11069 6502 11115 6554
rect 11115 6502 11125 6554
rect 11149 6502 11179 6554
rect 11179 6502 11191 6554
rect 11191 6502 11205 6554
rect 11229 6502 11243 6554
rect 11243 6502 11255 6554
rect 11255 6502 11285 6554
rect 11309 6502 11319 6554
rect 11319 6502 11365 6554
rect 11069 6500 11125 6502
rect 11149 6500 11205 6502
rect 11229 6500 11285 6502
rect 11309 6500 11365 6502
rect 11069 5466 11125 5468
rect 11149 5466 11205 5468
rect 11229 5466 11285 5468
rect 11309 5466 11365 5468
rect 11069 5414 11115 5466
rect 11115 5414 11125 5466
rect 11149 5414 11179 5466
rect 11179 5414 11191 5466
rect 11191 5414 11205 5466
rect 11229 5414 11243 5466
rect 11243 5414 11255 5466
rect 11255 5414 11285 5466
rect 11309 5414 11319 5466
rect 11319 5414 11365 5466
rect 11069 5412 11125 5414
rect 11149 5412 11205 5414
rect 11229 5412 11285 5414
rect 11309 5412 11365 5414
rect 11069 4378 11125 4380
rect 11149 4378 11205 4380
rect 11229 4378 11285 4380
rect 11309 4378 11365 4380
rect 11069 4326 11115 4378
rect 11115 4326 11125 4378
rect 11149 4326 11179 4378
rect 11179 4326 11191 4378
rect 11191 4326 11205 4378
rect 11229 4326 11243 4378
rect 11243 4326 11255 4378
rect 11255 4326 11285 4378
rect 11309 4326 11319 4378
rect 11319 4326 11365 4378
rect 11069 4324 11125 4326
rect 11149 4324 11205 4326
rect 11229 4324 11285 4326
rect 11309 4324 11365 4326
rect 11069 3290 11125 3292
rect 11149 3290 11205 3292
rect 11229 3290 11285 3292
rect 11309 3290 11365 3292
rect 11069 3238 11115 3290
rect 11115 3238 11125 3290
rect 11149 3238 11179 3290
rect 11179 3238 11191 3290
rect 11191 3238 11205 3290
rect 11229 3238 11243 3290
rect 11243 3238 11255 3290
rect 11255 3238 11285 3290
rect 11309 3238 11319 3290
rect 11319 3238 11365 3290
rect 11069 3236 11125 3238
rect 11149 3236 11205 3238
rect 11229 3236 11285 3238
rect 11309 3236 11365 3238
rect 14278 20848 14334 20884
rect 12622 15036 12624 15056
rect 12624 15036 12676 15056
rect 12676 15036 12678 15056
rect 12622 15000 12678 15036
rect 14462 18844 14464 18864
rect 14464 18844 14516 18864
rect 14516 18844 14518 18864
rect 14462 18808 14518 18844
rect 14646 18284 14702 18320
rect 14646 18264 14648 18284
rect 14648 18264 14700 18284
rect 14700 18264 14702 18284
rect 16711 25594 16767 25596
rect 16791 25594 16847 25596
rect 16871 25594 16927 25596
rect 16951 25594 17007 25596
rect 16711 25542 16757 25594
rect 16757 25542 16767 25594
rect 16791 25542 16821 25594
rect 16821 25542 16833 25594
rect 16833 25542 16847 25594
rect 16871 25542 16885 25594
rect 16885 25542 16897 25594
rect 16897 25542 16927 25594
rect 16951 25542 16961 25594
rect 16961 25542 17007 25594
rect 16711 25540 16767 25542
rect 16791 25540 16847 25542
rect 16871 25540 16927 25542
rect 16951 25540 17007 25542
rect 17371 26138 17427 26140
rect 17451 26138 17507 26140
rect 17531 26138 17587 26140
rect 17611 26138 17667 26140
rect 17371 26086 17417 26138
rect 17417 26086 17427 26138
rect 17451 26086 17481 26138
rect 17481 26086 17493 26138
rect 17493 26086 17507 26138
rect 17531 26086 17545 26138
rect 17545 26086 17557 26138
rect 17557 26086 17587 26138
rect 17611 26086 17621 26138
rect 17621 26086 17667 26138
rect 17371 26084 17427 26086
rect 17451 26084 17507 26086
rect 17531 26084 17587 26086
rect 17611 26084 17667 26086
rect 17371 25050 17427 25052
rect 17451 25050 17507 25052
rect 17531 25050 17587 25052
rect 17611 25050 17667 25052
rect 17371 24998 17417 25050
rect 17417 24998 17427 25050
rect 17451 24998 17481 25050
rect 17481 24998 17493 25050
rect 17493 24998 17507 25050
rect 17531 24998 17545 25050
rect 17545 24998 17557 25050
rect 17557 24998 17587 25050
rect 17611 24998 17621 25050
rect 17621 24998 17667 25050
rect 17371 24996 17427 24998
rect 17451 24996 17507 24998
rect 17531 24996 17587 24998
rect 17611 24996 17667 24998
rect 17130 24812 17186 24848
rect 17130 24792 17132 24812
rect 17132 24792 17184 24812
rect 17184 24792 17186 24812
rect 17774 24792 17830 24848
rect 16711 24506 16767 24508
rect 16791 24506 16847 24508
rect 16871 24506 16927 24508
rect 16951 24506 17007 24508
rect 16711 24454 16757 24506
rect 16757 24454 16767 24506
rect 16791 24454 16821 24506
rect 16821 24454 16833 24506
rect 16833 24454 16847 24506
rect 16871 24454 16885 24506
rect 16885 24454 16897 24506
rect 16897 24454 16927 24506
rect 16951 24454 16961 24506
rect 16961 24454 17007 24506
rect 16711 24452 16767 24454
rect 16791 24452 16847 24454
rect 16871 24452 16927 24454
rect 16951 24452 17007 24454
rect 17371 23962 17427 23964
rect 17451 23962 17507 23964
rect 17531 23962 17587 23964
rect 17611 23962 17667 23964
rect 17371 23910 17417 23962
rect 17417 23910 17427 23962
rect 17451 23910 17481 23962
rect 17481 23910 17493 23962
rect 17493 23910 17507 23962
rect 17531 23910 17545 23962
rect 17545 23910 17557 23962
rect 17557 23910 17587 23962
rect 17611 23910 17621 23962
rect 17621 23910 17667 23962
rect 17371 23908 17427 23910
rect 17451 23908 17507 23910
rect 17531 23908 17587 23910
rect 17611 23908 17667 23910
rect 16711 23418 16767 23420
rect 16791 23418 16847 23420
rect 16871 23418 16927 23420
rect 16951 23418 17007 23420
rect 16711 23366 16757 23418
rect 16757 23366 16767 23418
rect 16791 23366 16821 23418
rect 16821 23366 16833 23418
rect 16833 23366 16847 23418
rect 16871 23366 16885 23418
rect 16885 23366 16897 23418
rect 16897 23366 16927 23418
rect 16951 23366 16961 23418
rect 16961 23366 17007 23418
rect 16711 23364 16767 23366
rect 16791 23364 16847 23366
rect 16871 23364 16927 23366
rect 16951 23364 17007 23366
rect 17371 22874 17427 22876
rect 17451 22874 17507 22876
rect 17531 22874 17587 22876
rect 17611 22874 17667 22876
rect 17371 22822 17417 22874
rect 17417 22822 17427 22874
rect 17451 22822 17481 22874
rect 17481 22822 17493 22874
rect 17493 22822 17507 22874
rect 17531 22822 17545 22874
rect 17545 22822 17557 22874
rect 17557 22822 17587 22874
rect 17611 22822 17621 22874
rect 17621 22822 17667 22874
rect 17371 22820 17427 22822
rect 17451 22820 17507 22822
rect 17531 22820 17587 22822
rect 17611 22820 17667 22822
rect 15198 20460 15254 20496
rect 15198 20440 15200 20460
rect 15200 20440 15252 20460
rect 15252 20440 15254 20460
rect 13910 4564 13912 4584
rect 13912 4564 13964 4584
rect 13964 4564 13966 4584
rect 13910 4528 13966 4564
rect 11069 2202 11125 2204
rect 11149 2202 11205 2204
rect 11229 2202 11285 2204
rect 11309 2202 11365 2204
rect 11069 2150 11115 2202
rect 11115 2150 11125 2202
rect 11149 2150 11179 2202
rect 11179 2150 11191 2202
rect 11191 2150 11205 2202
rect 11229 2150 11243 2202
rect 11243 2150 11255 2202
rect 11255 2150 11285 2202
rect 11309 2150 11319 2202
rect 11319 2150 11365 2202
rect 11069 2148 11125 2150
rect 11149 2148 11205 2150
rect 11229 2148 11285 2150
rect 11309 2148 11365 2150
rect 16118 18128 16174 18184
rect 16711 22330 16767 22332
rect 16791 22330 16847 22332
rect 16871 22330 16927 22332
rect 16951 22330 17007 22332
rect 16711 22278 16757 22330
rect 16757 22278 16767 22330
rect 16791 22278 16821 22330
rect 16821 22278 16833 22330
rect 16833 22278 16847 22330
rect 16871 22278 16885 22330
rect 16885 22278 16897 22330
rect 16897 22278 16927 22330
rect 16951 22278 16961 22330
rect 16961 22278 17007 22330
rect 16711 22276 16767 22278
rect 16791 22276 16847 22278
rect 16871 22276 16927 22278
rect 16951 22276 17007 22278
rect 16711 21242 16767 21244
rect 16791 21242 16847 21244
rect 16871 21242 16927 21244
rect 16951 21242 17007 21244
rect 16711 21190 16757 21242
rect 16757 21190 16767 21242
rect 16791 21190 16821 21242
rect 16821 21190 16833 21242
rect 16833 21190 16847 21242
rect 16871 21190 16885 21242
rect 16885 21190 16897 21242
rect 16897 21190 16927 21242
rect 16951 21190 16961 21242
rect 16961 21190 17007 21242
rect 16711 21188 16767 21190
rect 16791 21188 16847 21190
rect 16871 21188 16927 21190
rect 16951 21188 17007 21190
rect 16711 20154 16767 20156
rect 16791 20154 16847 20156
rect 16871 20154 16927 20156
rect 16951 20154 17007 20156
rect 16711 20102 16757 20154
rect 16757 20102 16767 20154
rect 16791 20102 16821 20154
rect 16821 20102 16833 20154
rect 16833 20102 16847 20154
rect 16871 20102 16885 20154
rect 16885 20102 16897 20154
rect 16897 20102 16927 20154
rect 16951 20102 16961 20154
rect 16961 20102 17007 20154
rect 16711 20100 16767 20102
rect 16791 20100 16847 20102
rect 16871 20100 16927 20102
rect 16951 20100 17007 20102
rect 17371 21786 17427 21788
rect 17451 21786 17507 21788
rect 17531 21786 17587 21788
rect 17611 21786 17667 21788
rect 17371 21734 17417 21786
rect 17417 21734 17427 21786
rect 17451 21734 17481 21786
rect 17481 21734 17493 21786
rect 17493 21734 17507 21786
rect 17531 21734 17545 21786
rect 17545 21734 17557 21786
rect 17557 21734 17587 21786
rect 17611 21734 17621 21786
rect 17621 21734 17667 21786
rect 17371 21732 17427 21734
rect 17451 21732 17507 21734
rect 17531 21732 17587 21734
rect 17611 21732 17667 21734
rect 17371 20698 17427 20700
rect 17451 20698 17507 20700
rect 17531 20698 17587 20700
rect 17611 20698 17667 20700
rect 17371 20646 17417 20698
rect 17417 20646 17427 20698
rect 17451 20646 17481 20698
rect 17481 20646 17493 20698
rect 17493 20646 17507 20698
rect 17531 20646 17545 20698
rect 17545 20646 17557 20698
rect 17557 20646 17587 20698
rect 17611 20646 17621 20698
rect 17621 20646 17667 20698
rect 17371 20644 17427 20646
rect 17451 20644 17507 20646
rect 17531 20644 17587 20646
rect 17611 20644 17667 20646
rect 17130 19760 17186 19816
rect 19062 20848 19118 20904
rect 17371 19610 17427 19612
rect 17451 19610 17507 19612
rect 17531 19610 17587 19612
rect 17611 19610 17667 19612
rect 17371 19558 17417 19610
rect 17417 19558 17427 19610
rect 17451 19558 17481 19610
rect 17481 19558 17493 19610
rect 17493 19558 17507 19610
rect 17531 19558 17545 19610
rect 17545 19558 17557 19610
rect 17557 19558 17587 19610
rect 17611 19558 17621 19610
rect 17621 19558 17667 19610
rect 17371 19556 17427 19558
rect 17451 19556 17507 19558
rect 17531 19556 17587 19558
rect 17611 19556 17667 19558
rect 16711 19066 16767 19068
rect 16791 19066 16847 19068
rect 16871 19066 16927 19068
rect 16951 19066 17007 19068
rect 16711 19014 16757 19066
rect 16757 19014 16767 19066
rect 16791 19014 16821 19066
rect 16821 19014 16833 19066
rect 16833 19014 16847 19066
rect 16871 19014 16885 19066
rect 16885 19014 16897 19066
rect 16897 19014 16927 19066
rect 16951 19014 16961 19066
rect 16961 19014 17007 19066
rect 16711 19012 16767 19014
rect 16791 19012 16847 19014
rect 16871 19012 16927 19014
rect 16951 19012 17007 19014
rect 16394 18400 16450 18456
rect 16711 17978 16767 17980
rect 16791 17978 16847 17980
rect 16871 17978 16927 17980
rect 16951 17978 17007 17980
rect 16711 17926 16757 17978
rect 16757 17926 16767 17978
rect 16791 17926 16821 17978
rect 16821 17926 16833 17978
rect 16833 17926 16847 17978
rect 16871 17926 16885 17978
rect 16885 17926 16897 17978
rect 16897 17926 16927 17978
rect 16951 17926 16961 17978
rect 16961 17926 17007 17978
rect 16711 17924 16767 17926
rect 16791 17924 16847 17926
rect 16871 17924 16927 17926
rect 16951 17924 17007 17926
rect 17371 18522 17427 18524
rect 17451 18522 17507 18524
rect 17531 18522 17587 18524
rect 17611 18522 17667 18524
rect 17371 18470 17417 18522
rect 17417 18470 17427 18522
rect 17451 18470 17481 18522
rect 17481 18470 17493 18522
rect 17493 18470 17507 18522
rect 17531 18470 17545 18522
rect 17545 18470 17557 18522
rect 17557 18470 17587 18522
rect 17611 18470 17621 18522
rect 17621 18470 17667 18522
rect 17371 18468 17427 18470
rect 17451 18468 17507 18470
rect 17531 18468 17587 18470
rect 17611 18468 17667 18470
rect 17222 18400 17278 18456
rect 17406 18128 17462 18184
rect 17371 17434 17427 17436
rect 17451 17434 17507 17436
rect 17531 17434 17587 17436
rect 17611 17434 17667 17436
rect 17371 17382 17417 17434
rect 17417 17382 17427 17434
rect 17451 17382 17481 17434
rect 17481 17382 17493 17434
rect 17493 17382 17507 17434
rect 17531 17382 17545 17434
rect 17545 17382 17557 17434
rect 17557 17382 17587 17434
rect 17611 17382 17621 17434
rect 17621 17382 17667 17434
rect 17371 17380 17427 17382
rect 17451 17380 17507 17382
rect 17531 17380 17587 17382
rect 17611 17380 17667 17382
rect 16711 16890 16767 16892
rect 16791 16890 16847 16892
rect 16871 16890 16927 16892
rect 16951 16890 17007 16892
rect 16711 16838 16757 16890
rect 16757 16838 16767 16890
rect 16791 16838 16821 16890
rect 16821 16838 16833 16890
rect 16833 16838 16847 16890
rect 16871 16838 16885 16890
rect 16885 16838 16897 16890
rect 16897 16838 16927 16890
rect 16951 16838 16961 16890
rect 16961 16838 17007 16890
rect 16711 16836 16767 16838
rect 16791 16836 16847 16838
rect 16871 16836 16927 16838
rect 16951 16836 17007 16838
rect 17371 16346 17427 16348
rect 17451 16346 17507 16348
rect 17531 16346 17587 16348
rect 17611 16346 17667 16348
rect 17371 16294 17417 16346
rect 17417 16294 17427 16346
rect 17451 16294 17481 16346
rect 17481 16294 17493 16346
rect 17493 16294 17507 16346
rect 17531 16294 17545 16346
rect 17545 16294 17557 16346
rect 17557 16294 17587 16346
rect 17611 16294 17621 16346
rect 17621 16294 17667 16346
rect 17371 16292 17427 16294
rect 17451 16292 17507 16294
rect 17531 16292 17587 16294
rect 17611 16292 17667 16294
rect 16711 15802 16767 15804
rect 16791 15802 16847 15804
rect 16871 15802 16927 15804
rect 16951 15802 17007 15804
rect 16711 15750 16757 15802
rect 16757 15750 16767 15802
rect 16791 15750 16821 15802
rect 16821 15750 16833 15802
rect 16833 15750 16847 15802
rect 16871 15750 16885 15802
rect 16885 15750 16897 15802
rect 16897 15750 16927 15802
rect 16951 15750 16961 15802
rect 16961 15750 17007 15802
rect 16711 15748 16767 15750
rect 16791 15748 16847 15750
rect 16871 15748 16927 15750
rect 16951 15748 17007 15750
rect 16711 14714 16767 14716
rect 16791 14714 16847 14716
rect 16871 14714 16927 14716
rect 16951 14714 17007 14716
rect 16711 14662 16757 14714
rect 16757 14662 16767 14714
rect 16791 14662 16821 14714
rect 16821 14662 16833 14714
rect 16833 14662 16847 14714
rect 16871 14662 16885 14714
rect 16885 14662 16897 14714
rect 16897 14662 16927 14714
rect 16951 14662 16961 14714
rect 16961 14662 17007 14714
rect 16711 14660 16767 14662
rect 16791 14660 16847 14662
rect 16871 14660 16927 14662
rect 16951 14660 17007 14662
rect 23013 26682 23069 26684
rect 23093 26682 23149 26684
rect 23173 26682 23229 26684
rect 23253 26682 23309 26684
rect 23013 26630 23059 26682
rect 23059 26630 23069 26682
rect 23093 26630 23123 26682
rect 23123 26630 23135 26682
rect 23135 26630 23149 26682
rect 23173 26630 23187 26682
rect 23187 26630 23199 26682
rect 23199 26630 23229 26682
rect 23253 26630 23263 26682
rect 23263 26630 23309 26682
rect 23013 26628 23069 26630
rect 23093 26628 23149 26630
rect 23173 26628 23229 26630
rect 23253 26628 23309 26630
rect 23673 26138 23729 26140
rect 23753 26138 23809 26140
rect 23833 26138 23889 26140
rect 23913 26138 23969 26140
rect 23673 26086 23719 26138
rect 23719 26086 23729 26138
rect 23753 26086 23783 26138
rect 23783 26086 23795 26138
rect 23795 26086 23809 26138
rect 23833 26086 23847 26138
rect 23847 26086 23859 26138
rect 23859 26086 23889 26138
rect 23913 26086 23923 26138
rect 23923 26086 23969 26138
rect 23673 26084 23729 26086
rect 23753 26084 23809 26086
rect 23833 26084 23889 26086
rect 23913 26084 23969 26086
rect 20258 24112 20314 24168
rect 20074 23180 20130 23216
rect 20074 23160 20076 23180
rect 20076 23160 20128 23180
rect 20128 23160 20130 23180
rect 20350 23296 20406 23352
rect 19890 23044 19946 23080
rect 19890 23024 19892 23044
rect 19892 23024 19944 23044
rect 19944 23024 19946 23044
rect 20718 23316 20774 23352
rect 20718 23296 20720 23316
rect 20720 23296 20772 23316
rect 20772 23296 20774 23316
rect 20718 23180 20774 23216
rect 20718 23160 20720 23180
rect 20720 23160 20772 23180
rect 20772 23160 20774 23180
rect 21270 23024 21326 23080
rect 23013 25594 23069 25596
rect 23093 25594 23149 25596
rect 23173 25594 23229 25596
rect 23253 25594 23309 25596
rect 23013 25542 23059 25594
rect 23059 25542 23069 25594
rect 23093 25542 23123 25594
rect 23123 25542 23135 25594
rect 23135 25542 23149 25594
rect 23173 25542 23187 25594
rect 23187 25542 23199 25594
rect 23199 25542 23229 25594
rect 23253 25542 23263 25594
rect 23263 25542 23309 25594
rect 23013 25540 23069 25542
rect 23093 25540 23149 25542
rect 23173 25540 23229 25542
rect 23253 25540 23309 25542
rect 25778 25236 25780 25256
rect 25780 25236 25832 25256
rect 25832 25236 25834 25256
rect 19430 20848 19486 20904
rect 17371 15258 17427 15260
rect 17451 15258 17507 15260
rect 17531 15258 17587 15260
rect 17611 15258 17667 15260
rect 17371 15206 17417 15258
rect 17417 15206 17427 15258
rect 17451 15206 17481 15258
rect 17481 15206 17493 15258
rect 17493 15206 17507 15258
rect 17531 15206 17545 15258
rect 17545 15206 17557 15258
rect 17557 15206 17587 15258
rect 17611 15206 17621 15258
rect 17621 15206 17667 15258
rect 17371 15204 17427 15206
rect 17451 15204 17507 15206
rect 17531 15204 17587 15206
rect 17611 15204 17667 15206
rect 17371 14170 17427 14172
rect 17451 14170 17507 14172
rect 17531 14170 17587 14172
rect 17611 14170 17667 14172
rect 17371 14118 17417 14170
rect 17417 14118 17427 14170
rect 17451 14118 17481 14170
rect 17481 14118 17493 14170
rect 17493 14118 17507 14170
rect 17531 14118 17545 14170
rect 17545 14118 17557 14170
rect 17557 14118 17587 14170
rect 17611 14118 17621 14170
rect 17621 14118 17667 14170
rect 17371 14116 17427 14118
rect 17451 14116 17507 14118
rect 17531 14116 17587 14118
rect 17611 14116 17667 14118
rect 16711 13626 16767 13628
rect 16791 13626 16847 13628
rect 16871 13626 16927 13628
rect 16951 13626 17007 13628
rect 16711 13574 16757 13626
rect 16757 13574 16767 13626
rect 16791 13574 16821 13626
rect 16821 13574 16833 13626
rect 16833 13574 16847 13626
rect 16871 13574 16885 13626
rect 16885 13574 16897 13626
rect 16897 13574 16927 13626
rect 16951 13574 16961 13626
rect 16961 13574 17007 13626
rect 16711 13572 16767 13574
rect 16791 13572 16847 13574
rect 16871 13572 16927 13574
rect 16951 13572 17007 13574
rect 16711 12538 16767 12540
rect 16791 12538 16847 12540
rect 16871 12538 16927 12540
rect 16951 12538 17007 12540
rect 16711 12486 16757 12538
rect 16757 12486 16767 12538
rect 16791 12486 16821 12538
rect 16821 12486 16833 12538
rect 16833 12486 16847 12538
rect 16871 12486 16885 12538
rect 16885 12486 16897 12538
rect 16897 12486 16927 12538
rect 16951 12486 16961 12538
rect 16961 12486 17007 12538
rect 16711 12484 16767 12486
rect 16791 12484 16847 12486
rect 16871 12484 16927 12486
rect 16951 12484 17007 12486
rect 15106 9016 15162 9072
rect 17371 13082 17427 13084
rect 17451 13082 17507 13084
rect 17531 13082 17587 13084
rect 17611 13082 17667 13084
rect 17371 13030 17417 13082
rect 17417 13030 17427 13082
rect 17451 13030 17481 13082
rect 17481 13030 17493 13082
rect 17493 13030 17507 13082
rect 17531 13030 17545 13082
rect 17545 13030 17557 13082
rect 17557 13030 17587 13082
rect 17611 13030 17621 13082
rect 17621 13030 17667 13082
rect 17371 13028 17427 13030
rect 17451 13028 17507 13030
rect 17531 13028 17587 13030
rect 17611 13028 17667 13030
rect 16711 11450 16767 11452
rect 16791 11450 16847 11452
rect 16871 11450 16927 11452
rect 16951 11450 17007 11452
rect 16711 11398 16757 11450
rect 16757 11398 16767 11450
rect 16791 11398 16821 11450
rect 16821 11398 16833 11450
rect 16833 11398 16847 11450
rect 16871 11398 16885 11450
rect 16885 11398 16897 11450
rect 16897 11398 16927 11450
rect 16951 11398 16961 11450
rect 16961 11398 17007 11450
rect 16711 11396 16767 11398
rect 16791 11396 16847 11398
rect 16871 11396 16927 11398
rect 16951 11396 17007 11398
rect 16711 10362 16767 10364
rect 16791 10362 16847 10364
rect 16871 10362 16927 10364
rect 16951 10362 17007 10364
rect 16711 10310 16757 10362
rect 16757 10310 16767 10362
rect 16791 10310 16821 10362
rect 16821 10310 16833 10362
rect 16833 10310 16847 10362
rect 16871 10310 16885 10362
rect 16885 10310 16897 10362
rect 16897 10310 16927 10362
rect 16951 10310 16961 10362
rect 16961 10310 17007 10362
rect 16711 10308 16767 10310
rect 16791 10308 16847 10310
rect 16871 10308 16927 10310
rect 16951 10308 17007 10310
rect 16711 9274 16767 9276
rect 16791 9274 16847 9276
rect 16871 9274 16927 9276
rect 16951 9274 17007 9276
rect 16711 9222 16757 9274
rect 16757 9222 16767 9274
rect 16791 9222 16821 9274
rect 16821 9222 16833 9274
rect 16833 9222 16847 9274
rect 16871 9222 16885 9274
rect 16885 9222 16897 9274
rect 16897 9222 16927 9274
rect 16951 9222 16961 9274
rect 16961 9222 17007 9274
rect 16711 9220 16767 9222
rect 16791 9220 16847 9222
rect 16871 9220 16927 9222
rect 16951 9220 17007 9222
rect 17371 11994 17427 11996
rect 17451 11994 17507 11996
rect 17531 11994 17587 11996
rect 17611 11994 17667 11996
rect 17371 11942 17417 11994
rect 17417 11942 17427 11994
rect 17451 11942 17481 11994
rect 17481 11942 17493 11994
rect 17493 11942 17507 11994
rect 17531 11942 17545 11994
rect 17545 11942 17557 11994
rect 17557 11942 17587 11994
rect 17611 11942 17621 11994
rect 17621 11942 17667 11994
rect 17371 11940 17427 11942
rect 17451 11940 17507 11942
rect 17531 11940 17587 11942
rect 17611 11940 17667 11942
rect 17371 10906 17427 10908
rect 17451 10906 17507 10908
rect 17531 10906 17587 10908
rect 17611 10906 17667 10908
rect 17371 10854 17417 10906
rect 17417 10854 17427 10906
rect 17451 10854 17481 10906
rect 17481 10854 17493 10906
rect 17493 10854 17507 10906
rect 17531 10854 17545 10906
rect 17545 10854 17557 10906
rect 17557 10854 17587 10906
rect 17611 10854 17621 10906
rect 17621 10854 17667 10906
rect 17371 10852 17427 10854
rect 17451 10852 17507 10854
rect 17531 10852 17587 10854
rect 17611 10852 17667 10854
rect 17371 9818 17427 9820
rect 17451 9818 17507 9820
rect 17531 9818 17587 9820
rect 17611 9818 17667 9820
rect 17371 9766 17417 9818
rect 17417 9766 17427 9818
rect 17451 9766 17481 9818
rect 17481 9766 17493 9818
rect 17493 9766 17507 9818
rect 17531 9766 17545 9818
rect 17545 9766 17557 9818
rect 17557 9766 17587 9818
rect 17611 9766 17621 9818
rect 17621 9766 17667 9818
rect 17371 9764 17427 9766
rect 17451 9764 17507 9766
rect 17531 9764 17587 9766
rect 17611 9764 17667 9766
rect 20258 16632 20314 16688
rect 20718 16532 20720 16552
rect 20720 16532 20772 16552
rect 20772 16532 20774 16552
rect 20718 16496 20774 16532
rect 23013 24506 23069 24508
rect 23093 24506 23149 24508
rect 23173 24506 23229 24508
rect 23253 24506 23309 24508
rect 23013 24454 23059 24506
rect 23059 24454 23069 24506
rect 23093 24454 23123 24506
rect 23123 24454 23135 24506
rect 23135 24454 23149 24506
rect 23173 24454 23187 24506
rect 23187 24454 23199 24506
rect 23199 24454 23229 24506
rect 23253 24454 23263 24506
rect 23263 24454 23309 24506
rect 23013 24452 23069 24454
rect 23093 24452 23149 24454
rect 23173 24452 23229 24454
rect 23253 24452 23309 24454
rect 23110 24148 23112 24168
rect 23112 24148 23164 24168
rect 23164 24148 23166 24168
rect 23110 24112 23166 24148
rect 23673 25050 23729 25052
rect 23753 25050 23809 25052
rect 23833 25050 23889 25052
rect 23913 25050 23969 25052
rect 23673 24998 23719 25050
rect 23719 24998 23729 25050
rect 23753 24998 23783 25050
rect 23783 24998 23795 25050
rect 23795 24998 23809 25050
rect 23833 24998 23847 25050
rect 23847 24998 23859 25050
rect 23859 24998 23889 25050
rect 23913 24998 23923 25050
rect 23923 24998 23969 25050
rect 23673 24996 23729 24998
rect 23753 24996 23809 24998
rect 23833 24996 23889 24998
rect 23913 24996 23969 24998
rect 25778 25200 25834 25236
rect 23013 23418 23069 23420
rect 23093 23418 23149 23420
rect 23173 23418 23229 23420
rect 23253 23418 23309 23420
rect 23013 23366 23059 23418
rect 23059 23366 23069 23418
rect 23093 23366 23123 23418
rect 23123 23366 23135 23418
rect 23135 23366 23149 23418
rect 23173 23366 23187 23418
rect 23187 23366 23199 23418
rect 23199 23366 23229 23418
rect 23253 23366 23263 23418
rect 23263 23366 23309 23418
rect 23013 23364 23069 23366
rect 23093 23364 23149 23366
rect 23173 23364 23229 23366
rect 23253 23364 23309 23366
rect 23754 24132 23810 24168
rect 23754 24112 23756 24132
rect 23756 24112 23808 24132
rect 23808 24112 23810 24132
rect 23673 23962 23729 23964
rect 23753 23962 23809 23964
rect 23833 23962 23889 23964
rect 23913 23962 23969 23964
rect 23673 23910 23719 23962
rect 23719 23910 23729 23962
rect 23753 23910 23783 23962
rect 23783 23910 23795 23962
rect 23795 23910 23809 23962
rect 23833 23910 23847 23962
rect 23847 23910 23859 23962
rect 23859 23910 23889 23962
rect 23913 23910 23923 23962
rect 23923 23910 23969 23962
rect 23673 23908 23729 23910
rect 23753 23908 23809 23910
rect 23833 23908 23889 23910
rect 23913 23908 23969 23910
rect 23673 22874 23729 22876
rect 23753 22874 23809 22876
rect 23833 22874 23889 22876
rect 23913 22874 23969 22876
rect 23673 22822 23719 22874
rect 23719 22822 23729 22874
rect 23753 22822 23783 22874
rect 23783 22822 23795 22874
rect 23795 22822 23809 22874
rect 23833 22822 23847 22874
rect 23847 22822 23859 22874
rect 23859 22822 23889 22874
rect 23913 22822 23923 22874
rect 23923 22822 23969 22874
rect 23673 22820 23729 22822
rect 23753 22820 23809 22822
rect 23833 22820 23889 22822
rect 23913 22820 23969 22822
rect 23013 22330 23069 22332
rect 23093 22330 23149 22332
rect 23173 22330 23229 22332
rect 23253 22330 23309 22332
rect 23013 22278 23059 22330
rect 23059 22278 23069 22330
rect 23093 22278 23123 22330
rect 23123 22278 23135 22330
rect 23135 22278 23149 22330
rect 23173 22278 23187 22330
rect 23187 22278 23199 22330
rect 23199 22278 23229 22330
rect 23253 22278 23263 22330
rect 23263 22278 23309 22330
rect 23013 22276 23069 22278
rect 23093 22276 23149 22278
rect 23173 22276 23229 22278
rect 23253 22276 23309 22278
rect 23673 21786 23729 21788
rect 23753 21786 23809 21788
rect 23833 21786 23889 21788
rect 23913 21786 23969 21788
rect 23673 21734 23719 21786
rect 23719 21734 23729 21786
rect 23753 21734 23783 21786
rect 23783 21734 23795 21786
rect 23795 21734 23809 21786
rect 23833 21734 23847 21786
rect 23847 21734 23859 21786
rect 23859 21734 23889 21786
rect 23913 21734 23923 21786
rect 23923 21734 23969 21786
rect 23673 21732 23729 21734
rect 23753 21732 23809 21734
rect 23833 21732 23889 21734
rect 23913 21732 23969 21734
rect 23013 21242 23069 21244
rect 23093 21242 23149 21244
rect 23173 21242 23229 21244
rect 23253 21242 23309 21244
rect 23013 21190 23059 21242
rect 23059 21190 23069 21242
rect 23093 21190 23123 21242
rect 23123 21190 23135 21242
rect 23135 21190 23149 21242
rect 23173 21190 23187 21242
rect 23187 21190 23199 21242
rect 23199 21190 23229 21242
rect 23253 21190 23263 21242
rect 23263 21190 23309 21242
rect 23013 21188 23069 21190
rect 23093 21188 23149 21190
rect 23173 21188 23229 21190
rect 23253 21188 23309 21190
rect 23013 20154 23069 20156
rect 23093 20154 23149 20156
rect 23173 20154 23229 20156
rect 23253 20154 23309 20156
rect 23013 20102 23059 20154
rect 23059 20102 23069 20154
rect 23093 20102 23123 20154
rect 23123 20102 23135 20154
rect 23135 20102 23149 20154
rect 23173 20102 23187 20154
rect 23187 20102 23199 20154
rect 23199 20102 23229 20154
rect 23253 20102 23263 20154
rect 23263 20102 23309 20154
rect 23013 20100 23069 20102
rect 23093 20100 23149 20102
rect 23173 20100 23229 20102
rect 23253 20100 23309 20102
rect 23673 20698 23729 20700
rect 23753 20698 23809 20700
rect 23833 20698 23889 20700
rect 23913 20698 23969 20700
rect 23673 20646 23719 20698
rect 23719 20646 23729 20698
rect 23753 20646 23783 20698
rect 23783 20646 23795 20698
rect 23795 20646 23809 20698
rect 23833 20646 23847 20698
rect 23847 20646 23859 20698
rect 23859 20646 23889 20698
rect 23913 20646 23923 20698
rect 23923 20646 23969 20698
rect 23673 20644 23729 20646
rect 23753 20644 23809 20646
rect 23833 20644 23889 20646
rect 23913 20644 23969 20646
rect 23673 19610 23729 19612
rect 23753 19610 23809 19612
rect 23833 19610 23889 19612
rect 23913 19610 23969 19612
rect 23673 19558 23719 19610
rect 23719 19558 23729 19610
rect 23753 19558 23783 19610
rect 23783 19558 23795 19610
rect 23795 19558 23809 19610
rect 23833 19558 23847 19610
rect 23847 19558 23859 19610
rect 23859 19558 23889 19610
rect 23913 19558 23923 19610
rect 23923 19558 23969 19610
rect 23673 19556 23729 19558
rect 23753 19556 23809 19558
rect 23833 19556 23889 19558
rect 23913 19556 23969 19558
rect 23013 19066 23069 19068
rect 23093 19066 23149 19068
rect 23173 19066 23229 19068
rect 23253 19066 23309 19068
rect 23013 19014 23059 19066
rect 23059 19014 23069 19066
rect 23093 19014 23123 19066
rect 23123 19014 23135 19066
rect 23135 19014 23149 19066
rect 23173 19014 23187 19066
rect 23187 19014 23199 19066
rect 23199 19014 23229 19066
rect 23253 19014 23263 19066
rect 23263 19014 23309 19066
rect 23013 19012 23069 19014
rect 23093 19012 23149 19014
rect 23173 19012 23229 19014
rect 23253 19012 23309 19014
rect 22742 18808 22798 18864
rect 23013 17978 23069 17980
rect 23093 17978 23149 17980
rect 23173 17978 23229 17980
rect 23253 17978 23309 17980
rect 23013 17926 23059 17978
rect 23059 17926 23069 17978
rect 23093 17926 23123 17978
rect 23123 17926 23135 17978
rect 23135 17926 23149 17978
rect 23173 17926 23187 17978
rect 23187 17926 23199 17978
rect 23199 17926 23229 17978
rect 23253 17926 23263 17978
rect 23263 17926 23309 17978
rect 23013 17924 23069 17926
rect 23093 17924 23149 17926
rect 23173 17924 23229 17926
rect 23253 17924 23309 17926
rect 23673 18522 23729 18524
rect 23753 18522 23809 18524
rect 23833 18522 23889 18524
rect 23913 18522 23969 18524
rect 23673 18470 23719 18522
rect 23719 18470 23729 18522
rect 23753 18470 23783 18522
rect 23783 18470 23795 18522
rect 23795 18470 23809 18522
rect 23833 18470 23847 18522
rect 23847 18470 23859 18522
rect 23859 18470 23889 18522
rect 23913 18470 23923 18522
rect 23923 18470 23969 18522
rect 23673 18468 23729 18470
rect 23753 18468 23809 18470
rect 23833 18468 23889 18470
rect 23913 18468 23969 18470
rect 27066 23704 27122 23760
rect 25778 21120 25834 21176
rect 25226 18264 25282 18320
rect 21270 16532 21272 16552
rect 21272 16532 21324 16552
rect 21324 16532 21326 16552
rect 21270 16496 21326 16532
rect 23013 16890 23069 16892
rect 23093 16890 23149 16892
rect 23173 16890 23229 16892
rect 23253 16890 23309 16892
rect 23013 16838 23059 16890
rect 23059 16838 23069 16890
rect 23093 16838 23123 16890
rect 23123 16838 23135 16890
rect 23135 16838 23149 16890
rect 23173 16838 23187 16890
rect 23187 16838 23199 16890
rect 23199 16838 23229 16890
rect 23253 16838 23263 16890
rect 23263 16838 23309 16890
rect 23013 16836 23069 16838
rect 23093 16836 23149 16838
rect 23173 16836 23229 16838
rect 23253 16836 23309 16838
rect 23202 16668 23204 16688
rect 23204 16668 23256 16688
rect 23256 16668 23258 16688
rect 23202 16632 23258 16668
rect 23013 15802 23069 15804
rect 23093 15802 23149 15804
rect 23173 15802 23229 15804
rect 23253 15802 23309 15804
rect 23013 15750 23059 15802
rect 23059 15750 23069 15802
rect 23093 15750 23123 15802
rect 23123 15750 23135 15802
rect 23135 15750 23149 15802
rect 23173 15750 23187 15802
rect 23187 15750 23199 15802
rect 23199 15750 23229 15802
rect 23253 15750 23263 15802
rect 23263 15750 23309 15802
rect 23013 15748 23069 15750
rect 23093 15748 23149 15750
rect 23173 15748 23229 15750
rect 23253 15748 23309 15750
rect 23673 17434 23729 17436
rect 23753 17434 23809 17436
rect 23833 17434 23889 17436
rect 23913 17434 23969 17436
rect 23673 17382 23719 17434
rect 23719 17382 23729 17434
rect 23753 17382 23783 17434
rect 23783 17382 23795 17434
rect 23795 17382 23809 17434
rect 23833 17382 23847 17434
rect 23847 17382 23859 17434
rect 23859 17382 23889 17434
rect 23913 17382 23923 17434
rect 23923 17382 23969 17434
rect 23673 17380 23729 17382
rect 23753 17380 23809 17382
rect 23833 17380 23889 17382
rect 23913 17380 23969 17382
rect 23673 16346 23729 16348
rect 23753 16346 23809 16348
rect 23833 16346 23889 16348
rect 23913 16346 23969 16348
rect 23673 16294 23719 16346
rect 23719 16294 23729 16346
rect 23753 16294 23783 16346
rect 23783 16294 23795 16346
rect 23795 16294 23809 16346
rect 23833 16294 23847 16346
rect 23847 16294 23859 16346
rect 23859 16294 23889 16346
rect 23913 16294 23923 16346
rect 23923 16294 23969 16346
rect 23673 16292 23729 16294
rect 23753 16292 23809 16294
rect 23833 16292 23889 16294
rect 23913 16292 23969 16294
rect 23673 15258 23729 15260
rect 23753 15258 23809 15260
rect 23833 15258 23889 15260
rect 23913 15258 23969 15260
rect 23673 15206 23719 15258
rect 23719 15206 23729 15258
rect 23753 15206 23783 15258
rect 23783 15206 23795 15258
rect 23795 15206 23809 15258
rect 23833 15206 23847 15258
rect 23847 15206 23859 15258
rect 23859 15206 23889 15258
rect 23913 15206 23923 15258
rect 23923 15206 23969 15258
rect 23673 15204 23729 15206
rect 23753 15204 23809 15206
rect 23833 15204 23889 15206
rect 23913 15204 23969 15206
rect 23013 14714 23069 14716
rect 23093 14714 23149 14716
rect 23173 14714 23229 14716
rect 23253 14714 23309 14716
rect 23013 14662 23059 14714
rect 23059 14662 23069 14714
rect 23093 14662 23123 14714
rect 23123 14662 23135 14714
rect 23135 14662 23149 14714
rect 23173 14662 23187 14714
rect 23187 14662 23199 14714
rect 23199 14662 23229 14714
rect 23253 14662 23263 14714
rect 23263 14662 23309 14714
rect 23013 14660 23069 14662
rect 23093 14660 23149 14662
rect 23173 14660 23229 14662
rect 23253 14660 23309 14662
rect 23673 14170 23729 14172
rect 23753 14170 23809 14172
rect 23833 14170 23889 14172
rect 23913 14170 23969 14172
rect 23673 14118 23719 14170
rect 23719 14118 23729 14170
rect 23753 14118 23783 14170
rect 23783 14118 23795 14170
rect 23795 14118 23809 14170
rect 23833 14118 23847 14170
rect 23847 14118 23859 14170
rect 23859 14118 23889 14170
rect 23913 14118 23923 14170
rect 23923 14118 23969 14170
rect 23673 14116 23729 14118
rect 23753 14116 23809 14118
rect 23833 14116 23889 14118
rect 23913 14116 23969 14118
rect 23013 13626 23069 13628
rect 23093 13626 23149 13628
rect 23173 13626 23229 13628
rect 23253 13626 23309 13628
rect 23013 13574 23059 13626
rect 23059 13574 23069 13626
rect 23093 13574 23123 13626
rect 23123 13574 23135 13626
rect 23135 13574 23149 13626
rect 23173 13574 23187 13626
rect 23187 13574 23199 13626
rect 23199 13574 23229 13626
rect 23253 13574 23263 13626
rect 23263 13574 23309 13626
rect 23013 13572 23069 13574
rect 23093 13572 23149 13574
rect 23173 13572 23229 13574
rect 23253 13572 23309 13574
rect 16711 8186 16767 8188
rect 16791 8186 16847 8188
rect 16871 8186 16927 8188
rect 16951 8186 17007 8188
rect 16711 8134 16757 8186
rect 16757 8134 16767 8186
rect 16791 8134 16821 8186
rect 16821 8134 16833 8186
rect 16833 8134 16847 8186
rect 16871 8134 16885 8186
rect 16885 8134 16897 8186
rect 16897 8134 16927 8186
rect 16951 8134 16961 8186
rect 16961 8134 17007 8186
rect 16711 8132 16767 8134
rect 16791 8132 16847 8134
rect 16871 8132 16927 8134
rect 16951 8132 17007 8134
rect 15290 4564 15292 4584
rect 15292 4564 15344 4584
rect 15344 4564 15346 4584
rect 15290 4528 15346 4564
rect 16711 7098 16767 7100
rect 16791 7098 16847 7100
rect 16871 7098 16927 7100
rect 16951 7098 17007 7100
rect 16711 7046 16757 7098
rect 16757 7046 16767 7098
rect 16791 7046 16821 7098
rect 16821 7046 16833 7098
rect 16833 7046 16847 7098
rect 16871 7046 16885 7098
rect 16885 7046 16897 7098
rect 16897 7046 16927 7098
rect 16951 7046 16961 7098
rect 16961 7046 17007 7098
rect 16711 7044 16767 7046
rect 16791 7044 16847 7046
rect 16871 7044 16927 7046
rect 16951 7044 17007 7046
rect 17371 8730 17427 8732
rect 17451 8730 17507 8732
rect 17531 8730 17587 8732
rect 17611 8730 17667 8732
rect 17371 8678 17417 8730
rect 17417 8678 17427 8730
rect 17451 8678 17481 8730
rect 17481 8678 17493 8730
rect 17493 8678 17507 8730
rect 17531 8678 17545 8730
rect 17545 8678 17557 8730
rect 17557 8678 17587 8730
rect 17611 8678 17621 8730
rect 17621 8678 17667 8730
rect 17371 8676 17427 8678
rect 17451 8676 17507 8678
rect 17531 8676 17587 8678
rect 17611 8676 17667 8678
rect 17371 7642 17427 7644
rect 17451 7642 17507 7644
rect 17531 7642 17587 7644
rect 17611 7642 17667 7644
rect 17371 7590 17417 7642
rect 17417 7590 17427 7642
rect 17451 7590 17481 7642
rect 17481 7590 17493 7642
rect 17493 7590 17507 7642
rect 17531 7590 17545 7642
rect 17545 7590 17557 7642
rect 17557 7590 17587 7642
rect 17611 7590 17621 7642
rect 17621 7590 17667 7642
rect 17371 7588 17427 7590
rect 17451 7588 17507 7590
rect 17531 7588 17587 7590
rect 17611 7588 17667 7590
rect 20718 11736 20774 11792
rect 17371 6554 17427 6556
rect 17451 6554 17507 6556
rect 17531 6554 17587 6556
rect 17611 6554 17667 6556
rect 17371 6502 17417 6554
rect 17417 6502 17427 6554
rect 17451 6502 17481 6554
rect 17481 6502 17493 6554
rect 17493 6502 17507 6554
rect 17531 6502 17545 6554
rect 17545 6502 17557 6554
rect 17557 6502 17587 6554
rect 17611 6502 17621 6554
rect 17621 6502 17667 6554
rect 17371 6500 17427 6502
rect 17451 6500 17507 6502
rect 17531 6500 17587 6502
rect 17611 6500 17667 6502
rect 16711 6010 16767 6012
rect 16791 6010 16847 6012
rect 16871 6010 16927 6012
rect 16951 6010 17007 6012
rect 16711 5958 16757 6010
rect 16757 5958 16767 6010
rect 16791 5958 16821 6010
rect 16821 5958 16833 6010
rect 16833 5958 16847 6010
rect 16871 5958 16885 6010
rect 16885 5958 16897 6010
rect 16897 5958 16927 6010
rect 16951 5958 16961 6010
rect 16961 5958 17007 6010
rect 16711 5956 16767 5958
rect 16791 5956 16847 5958
rect 16871 5956 16927 5958
rect 16951 5956 17007 5958
rect 17371 5466 17427 5468
rect 17451 5466 17507 5468
rect 17531 5466 17587 5468
rect 17611 5466 17667 5468
rect 17371 5414 17417 5466
rect 17417 5414 17427 5466
rect 17451 5414 17481 5466
rect 17481 5414 17493 5466
rect 17493 5414 17507 5466
rect 17531 5414 17545 5466
rect 17545 5414 17557 5466
rect 17557 5414 17587 5466
rect 17611 5414 17621 5466
rect 17621 5414 17667 5466
rect 17371 5412 17427 5414
rect 17451 5412 17507 5414
rect 17531 5412 17587 5414
rect 17611 5412 17667 5414
rect 17130 5244 17132 5264
rect 17132 5244 17184 5264
rect 17184 5244 17186 5264
rect 17130 5208 17186 5244
rect 17406 5228 17462 5264
rect 17406 5208 17408 5228
rect 17408 5208 17460 5228
rect 17460 5208 17462 5228
rect 16711 4922 16767 4924
rect 16791 4922 16847 4924
rect 16871 4922 16927 4924
rect 16951 4922 17007 4924
rect 16711 4870 16757 4922
rect 16757 4870 16767 4922
rect 16791 4870 16821 4922
rect 16821 4870 16833 4922
rect 16833 4870 16847 4922
rect 16871 4870 16885 4922
rect 16885 4870 16897 4922
rect 16897 4870 16927 4922
rect 16951 4870 16961 4922
rect 16961 4870 17007 4922
rect 16711 4868 16767 4870
rect 16791 4868 16847 4870
rect 16871 4868 16927 4870
rect 16951 4868 17007 4870
rect 17371 4378 17427 4380
rect 17451 4378 17507 4380
rect 17531 4378 17587 4380
rect 17611 4378 17667 4380
rect 17371 4326 17417 4378
rect 17417 4326 17427 4378
rect 17451 4326 17481 4378
rect 17481 4326 17493 4378
rect 17493 4326 17507 4378
rect 17531 4326 17545 4378
rect 17545 4326 17557 4378
rect 17557 4326 17587 4378
rect 17611 4326 17621 4378
rect 17621 4326 17667 4378
rect 17371 4324 17427 4326
rect 17451 4324 17507 4326
rect 17531 4324 17587 4326
rect 17611 4324 17667 4326
rect 16711 3834 16767 3836
rect 16791 3834 16847 3836
rect 16871 3834 16927 3836
rect 16951 3834 17007 3836
rect 16711 3782 16757 3834
rect 16757 3782 16767 3834
rect 16791 3782 16821 3834
rect 16821 3782 16833 3834
rect 16833 3782 16847 3834
rect 16871 3782 16885 3834
rect 16885 3782 16897 3834
rect 16897 3782 16927 3834
rect 16951 3782 16961 3834
rect 16961 3782 17007 3834
rect 16711 3780 16767 3782
rect 16791 3780 16847 3782
rect 16871 3780 16927 3782
rect 16951 3780 17007 3782
rect 16711 2746 16767 2748
rect 16791 2746 16847 2748
rect 16871 2746 16927 2748
rect 16951 2746 17007 2748
rect 16711 2694 16757 2746
rect 16757 2694 16767 2746
rect 16791 2694 16821 2746
rect 16821 2694 16833 2746
rect 16833 2694 16847 2746
rect 16871 2694 16885 2746
rect 16885 2694 16897 2746
rect 16897 2694 16927 2746
rect 16951 2694 16961 2746
rect 16961 2694 17007 2746
rect 16711 2692 16767 2694
rect 16791 2692 16847 2694
rect 16871 2692 16927 2694
rect 16951 2692 17007 2694
rect 17371 3290 17427 3292
rect 17451 3290 17507 3292
rect 17531 3290 17587 3292
rect 17611 3290 17667 3292
rect 17371 3238 17417 3290
rect 17417 3238 17427 3290
rect 17451 3238 17481 3290
rect 17481 3238 17493 3290
rect 17493 3238 17507 3290
rect 17531 3238 17545 3290
rect 17545 3238 17557 3290
rect 17557 3238 17587 3290
rect 17611 3238 17621 3290
rect 17621 3238 17667 3290
rect 17371 3236 17427 3238
rect 17451 3236 17507 3238
rect 17531 3236 17587 3238
rect 17611 3236 17667 3238
rect 18786 9016 18842 9072
rect 19338 6180 19394 6216
rect 19338 6160 19340 6180
rect 19340 6160 19392 6180
rect 19392 6160 19394 6180
rect 23673 13082 23729 13084
rect 23753 13082 23809 13084
rect 23833 13082 23889 13084
rect 23913 13082 23969 13084
rect 23673 13030 23719 13082
rect 23719 13030 23729 13082
rect 23753 13030 23783 13082
rect 23783 13030 23795 13082
rect 23795 13030 23809 13082
rect 23833 13030 23847 13082
rect 23847 13030 23859 13082
rect 23859 13030 23889 13082
rect 23913 13030 23923 13082
rect 23923 13030 23969 13082
rect 23673 13028 23729 13030
rect 23753 13028 23809 13030
rect 23833 13028 23889 13030
rect 23913 13028 23969 13030
rect 23013 12538 23069 12540
rect 23093 12538 23149 12540
rect 23173 12538 23229 12540
rect 23253 12538 23309 12540
rect 23013 12486 23059 12538
rect 23059 12486 23069 12538
rect 23093 12486 23123 12538
rect 23123 12486 23135 12538
rect 23135 12486 23149 12538
rect 23173 12486 23187 12538
rect 23187 12486 23199 12538
rect 23199 12486 23229 12538
rect 23253 12486 23263 12538
rect 23263 12486 23309 12538
rect 23013 12484 23069 12486
rect 23093 12484 23149 12486
rect 23173 12484 23229 12486
rect 23253 12484 23309 12486
rect 23673 11994 23729 11996
rect 23753 11994 23809 11996
rect 23833 11994 23889 11996
rect 23913 11994 23969 11996
rect 23673 11942 23719 11994
rect 23719 11942 23729 11994
rect 23753 11942 23783 11994
rect 23783 11942 23795 11994
rect 23795 11942 23809 11994
rect 23833 11942 23847 11994
rect 23847 11942 23859 11994
rect 23859 11942 23889 11994
rect 23913 11942 23923 11994
rect 23923 11942 23969 11994
rect 23673 11940 23729 11942
rect 23753 11940 23809 11942
rect 23833 11940 23889 11942
rect 23913 11940 23969 11942
rect 23110 11756 23166 11792
rect 23110 11736 23112 11756
rect 23112 11736 23164 11756
rect 23164 11736 23166 11756
rect 23013 11450 23069 11452
rect 23093 11450 23149 11452
rect 23173 11450 23229 11452
rect 23253 11450 23309 11452
rect 23013 11398 23059 11450
rect 23059 11398 23069 11450
rect 23093 11398 23123 11450
rect 23123 11398 23135 11450
rect 23135 11398 23149 11450
rect 23173 11398 23187 11450
rect 23187 11398 23199 11450
rect 23199 11398 23229 11450
rect 23253 11398 23263 11450
rect 23263 11398 23309 11450
rect 23013 11396 23069 11398
rect 23093 11396 23149 11398
rect 23173 11396 23229 11398
rect 23253 11396 23309 11398
rect 23013 10362 23069 10364
rect 23093 10362 23149 10364
rect 23173 10362 23229 10364
rect 23253 10362 23309 10364
rect 23013 10310 23059 10362
rect 23059 10310 23069 10362
rect 23093 10310 23123 10362
rect 23123 10310 23135 10362
rect 23135 10310 23149 10362
rect 23173 10310 23187 10362
rect 23187 10310 23199 10362
rect 23199 10310 23229 10362
rect 23253 10310 23263 10362
rect 23263 10310 23309 10362
rect 23013 10308 23069 10310
rect 23093 10308 23149 10310
rect 23173 10308 23229 10310
rect 23253 10308 23309 10310
rect 23013 9274 23069 9276
rect 23093 9274 23149 9276
rect 23173 9274 23229 9276
rect 23253 9274 23309 9276
rect 23013 9222 23059 9274
rect 23059 9222 23069 9274
rect 23093 9222 23123 9274
rect 23123 9222 23135 9274
rect 23135 9222 23149 9274
rect 23173 9222 23187 9274
rect 23187 9222 23199 9274
rect 23199 9222 23229 9274
rect 23253 9222 23263 9274
rect 23263 9222 23309 9274
rect 23013 9220 23069 9222
rect 23093 9220 23149 9222
rect 23173 9220 23229 9222
rect 23253 9220 23309 9222
rect 23673 10906 23729 10908
rect 23753 10906 23809 10908
rect 23833 10906 23889 10908
rect 23913 10906 23969 10908
rect 23673 10854 23719 10906
rect 23719 10854 23729 10906
rect 23753 10854 23783 10906
rect 23783 10854 23795 10906
rect 23795 10854 23809 10906
rect 23833 10854 23847 10906
rect 23847 10854 23859 10906
rect 23859 10854 23889 10906
rect 23913 10854 23923 10906
rect 23923 10854 23969 10906
rect 23673 10852 23729 10854
rect 23753 10852 23809 10854
rect 23833 10852 23889 10854
rect 23913 10852 23969 10854
rect 23673 9818 23729 9820
rect 23753 9818 23809 9820
rect 23833 9818 23889 9820
rect 23913 9818 23969 9820
rect 23673 9766 23719 9818
rect 23719 9766 23729 9818
rect 23753 9766 23783 9818
rect 23783 9766 23795 9818
rect 23795 9766 23809 9818
rect 23833 9766 23847 9818
rect 23847 9766 23859 9818
rect 23859 9766 23889 9818
rect 23913 9766 23923 9818
rect 23923 9766 23969 9818
rect 23673 9764 23729 9766
rect 23753 9764 23809 9766
rect 23833 9764 23889 9766
rect 23913 9764 23969 9766
rect 23673 8730 23729 8732
rect 23753 8730 23809 8732
rect 23833 8730 23889 8732
rect 23913 8730 23969 8732
rect 23673 8678 23719 8730
rect 23719 8678 23729 8730
rect 23753 8678 23783 8730
rect 23783 8678 23795 8730
rect 23795 8678 23809 8730
rect 23833 8678 23847 8730
rect 23847 8678 23859 8730
rect 23859 8678 23889 8730
rect 23913 8678 23923 8730
rect 23923 8678 23969 8730
rect 23673 8676 23729 8678
rect 23753 8676 23809 8678
rect 23833 8676 23889 8678
rect 23913 8676 23969 8678
rect 23013 8186 23069 8188
rect 23093 8186 23149 8188
rect 23173 8186 23229 8188
rect 23253 8186 23309 8188
rect 23013 8134 23059 8186
rect 23059 8134 23069 8186
rect 23093 8134 23123 8186
rect 23123 8134 23135 8186
rect 23135 8134 23149 8186
rect 23173 8134 23187 8186
rect 23187 8134 23199 8186
rect 23199 8134 23229 8186
rect 23253 8134 23263 8186
rect 23263 8134 23309 8186
rect 23013 8132 23069 8134
rect 23093 8132 23149 8134
rect 23173 8132 23229 8134
rect 23253 8132 23309 8134
rect 23673 7642 23729 7644
rect 23753 7642 23809 7644
rect 23833 7642 23889 7644
rect 23913 7642 23969 7644
rect 23673 7590 23719 7642
rect 23719 7590 23729 7642
rect 23753 7590 23783 7642
rect 23783 7590 23795 7642
rect 23795 7590 23809 7642
rect 23833 7590 23847 7642
rect 23847 7590 23859 7642
rect 23859 7590 23889 7642
rect 23913 7590 23923 7642
rect 23923 7590 23969 7642
rect 23673 7588 23729 7590
rect 23753 7588 23809 7590
rect 23833 7588 23889 7590
rect 23913 7588 23969 7590
rect 19706 6316 19762 6352
rect 19706 6296 19708 6316
rect 19708 6296 19760 6316
rect 19760 6296 19762 6316
rect 19706 6060 19708 6080
rect 19708 6060 19760 6080
rect 19760 6060 19762 6080
rect 19706 6024 19762 6060
rect 20350 6196 20352 6216
rect 20352 6196 20404 6216
rect 20404 6196 20406 6216
rect 20350 6160 20406 6196
rect 20166 5616 20222 5672
rect 20810 6296 20866 6352
rect 20534 6024 20590 6080
rect 23013 7098 23069 7100
rect 23093 7098 23149 7100
rect 23173 7098 23229 7100
rect 23253 7098 23309 7100
rect 23013 7046 23059 7098
rect 23059 7046 23069 7098
rect 23093 7046 23123 7098
rect 23123 7046 23135 7098
rect 23135 7046 23149 7098
rect 23173 7046 23187 7098
rect 23187 7046 23199 7098
rect 23199 7046 23229 7098
rect 23253 7046 23263 7098
rect 23263 7046 23309 7098
rect 23013 7044 23069 7046
rect 23093 7044 23149 7046
rect 23173 7044 23229 7046
rect 23253 7044 23309 7046
rect 25870 17060 25926 17096
rect 25870 17040 25872 17060
rect 25872 17040 25924 17060
rect 25924 17040 25926 17060
rect 25778 12960 25834 13016
rect 25870 8200 25926 8256
rect 22374 6060 22376 6080
rect 22376 6060 22428 6080
rect 22428 6060 22430 6080
rect 22374 6024 22430 6060
rect 22558 5616 22614 5672
rect 23013 6010 23069 6012
rect 23093 6010 23149 6012
rect 23173 6010 23229 6012
rect 23253 6010 23309 6012
rect 23013 5958 23059 6010
rect 23059 5958 23069 6010
rect 23093 5958 23123 6010
rect 23123 5958 23135 6010
rect 23135 5958 23149 6010
rect 23173 5958 23187 6010
rect 23187 5958 23199 6010
rect 23199 5958 23229 6010
rect 23253 5958 23263 6010
rect 23263 5958 23309 6010
rect 23013 5956 23069 5958
rect 23093 5956 23149 5958
rect 23173 5956 23229 5958
rect 23253 5956 23309 5958
rect 23673 6554 23729 6556
rect 23753 6554 23809 6556
rect 23833 6554 23889 6556
rect 23913 6554 23969 6556
rect 23673 6502 23719 6554
rect 23719 6502 23729 6554
rect 23753 6502 23783 6554
rect 23783 6502 23795 6554
rect 23795 6502 23809 6554
rect 23833 6502 23847 6554
rect 23847 6502 23859 6554
rect 23859 6502 23889 6554
rect 23913 6502 23923 6554
rect 23923 6502 23969 6554
rect 23673 6500 23729 6502
rect 23753 6500 23809 6502
rect 23833 6500 23889 6502
rect 23913 6500 23969 6502
rect 23673 5466 23729 5468
rect 23753 5466 23809 5468
rect 23833 5466 23889 5468
rect 23913 5466 23969 5468
rect 23673 5414 23719 5466
rect 23719 5414 23729 5466
rect 23753 5414 23783 5466
rect 23783 5414 23795 5466
rect 23795 5414 23809 5466
rect 23833 5414 23847 5466
rect 23847 5414 23859 5466
rect 23859 5414 23889 5466
rect 23913 5414 23923 5466
rect 23923 5414 23969 5466
rect 23673 5412 23729 5414
rect 23753 5412 23809 5414
rect 23833 5412 23889 5414
rect 23913 5412 23969 5414
rect 23013 4922 23069 4924
rect 23093 4922 23149 4924
rect 23173 4922 23229 4924
rect 23253 4922 23309 4924
rect 23013 4870 23059 4922
rect 23059 4870 23069 4922
rect 23093 4870 23123 4922
rect 23123 4870 23135 4922
rect 23135 4870 23149 4922
rect 23173 4870 23187 4922
rect 23187 4870 23199 4922
rect 23199 4870 23229 4922
rect 23253 4870 23263 4922
rect 23263 4870 23309 4922
rect 23013 4868 23069 4870
rect 23093 4868 23149 4870
rect 23173 4868 23229 4870
rect 23253 4868 23309 4870
rect 23673 4378 23729 4380
rect 23753 4378 23809 4380
rect 23833 4378 23889 4380
rect 23913 4378 23969 4380
rect 23673 4326 23719 4378
rect 23719 4326 23729 4378
rect 23753 4326 23783 4378
rect 23783 4326 23795 4378
rect 23795 4326 23809 4378
rect 23833 4326 23847 4378
rect 23847 4326 23859 4378
rect 23859 4326 23889 4378
rect 23913 4326 23923 4378
rect 23923 4326 23969 4378
rect 23673 4324 23729 4326
rect 23753 4324 23809 4326
rect 23833 4324 23889 4326
rect 23913 4324 23969 4326
rect 23013 3834 23069 3836
rect 23093 3834 23149 3836
rect 23173 3834 23229 3836
rect 23253 3834 23309 3836
rect 23013 3782 23059 3834
rect 23059 3782 23069 3834
rect 23093 3782 23123 3834
rect 23123 3782 23135 3834
rect 23135 3782 23149 3834
rect 23173 3782 23187 3834
rect 23187 3782 23199 3834
rect 23199 3782 23229 3834
rect 23253 3782 23263 3834
rect 23263 3782 23309 3834
rect 23013 3780 23069 3782
rect 23093 3780 23149 3782
rect 23173 3780 23229 3782
rect 23253 3780 23309 3782
rect 25778 4120 25834 4176
rect 23013 2746 23069 2748
rect 23093 2746 23149 2748
rect 23173 2746 23229 2748
rect 23253 2746 23309 2748
rect 23013 2694 23059 2746
rect 23059 2694 23069 2746
rect 23093 2694 23123 2746
rect 23123 2694 23135 2746
rect 23135 2694 23149 2746
rect 23173 2694 23187 2746
rect 23187 2694 23199 2746
rect 23199 2694 23229 2746
rect 23253 2694 23263 2746
rect 23263 2694 23309 2746
rect 23013 2692 23069 2694
rect 23093 2692 23149 2694
rect 23173 2692 23229 2694
rect 23253 2692 23309 2694
rect 23673 3290 23729 3292
rect 23753 3290 23809 3292
rect 23833 3290 23889 3292
rect 23913 3290 23969 3292
rect 23673 3238 23719 3290
rect 23719 3238 23729 3290
rect 23753 3238 23783 3290
rect 23783 3238 23795 3290
rect 23795 3238 23809 3290
rect 23833 3238 23847 3290
rect 23847 3238 23859 3290
rect 23859 3238 23889 3290
rect 23913 3238 23923 3290
rect 23923 3238 23969 3290
rect 23673 3236 23729 3238
rect 23753 3236 23809 3238
rect 23833 3236 23889 3238
rect 23913 3236 23969 3238
rect 17371 2202 17427 2204
rect 17451 2202 17507 2204
rect 17531 2202 17587 2204
rect 17611 2202 17667 2204
rect 17371 2150 17417 2202
rect 17417 2150 17427 2202
rect 17451 2150 17481 2202
rect 17481 2150 17493 2202
rect 17493 2150 17507 2202
rect 17531 2150 17545 2202
rect 17545 2150 17557 2202
rect 17557 2150 17587 2202
rect 17611 2150 17621 2202
rect 17621 2150 17667 2202
rect 17371 2148 17427 2150
rect 17451 2148 17507 2150
rect 17531 2148 17587 2150
rect 17611 2148 17667 2150
rect 23673 2202 23729 2204
rect 23753 2202 23809 2204
rect 23833 2202 23889 2204
rect 23913 2202 23969 2204
rect 23673 2150 23719 2202
rect 23719 2150 23729 2202
rect 23753 2150 23783 2202
rect 23783 2150 23795 2202
rect 23795 2150 23809 2202
rect 23833 2150 23847 2202
rect 23847 2150 23859 2202
rect 23859 2150 23889 2202
rect 23913 2150 23923 2202
rect 23923 2150 23969 2202
rect 23673 2148 23729 2150
rect 23753 2148 23809 2150
rect 23833 2148 23889 2150
rect 23913 2148 23969 2150
rect 24766 40 24822 96
<< metal3 >>
rect 0 29338 800 29368
rect 1393 29338 1459 29341
rect 0 29336 1459 29338
rect 0 29280 1398 29336
rect 1454 29280 1459 29336
rect 0 29278 1459 29280
rect 0 29248 800 29278
rect 1393 29275 1459 29278
rect 4757 27232 5073 27233
rect 4757 27168 4763 27232
rect 4827 27168 4843 27232
rect 4907 27168 4923 27232
rect 4987 27168 5003 27232
rect 5067 27168 5073 27232
rect 4757 27167 5073 27168
rect 11059 27232 11375 27233
rect 11059 27168 11065 27232
rect 11129 27168 11145 27232
rect 11209 27168 11225 27232
rect 11289 27168 11305 27232
rect 11369 27168 11375 27232
rect 11059 27167 11375 27168
rect 17361 27232 17677 27233
rect 17361 27168 17367 27232
rect 17431 27168 17447 27232
rect 17511 27168 17527 27232
rect 17591 27168 17607 27232
rect 17671 27168 17677 27232
rect 17361 27167 17677 27168
rect 23663 27232 23979 27233
rect 23663 27168 23669 27232
rect 23733 27168 23749 27232
rect 23813 27168 23829 27232
rect 23893 27168 23909 27232
rect 23973 27168 23979 27232
rect 23663 27167 23979 27168
rect 4097 26688 4413 26689
rect 4097 26624 4103 26688
rect 4167 26624 4183 26688
rect 4247 26624 4263 26688
rect 4327 26624 4343 26688
rect 4407 26624 4413 26688
rect 4097 26623 4413 26624
rect 10399 26688 10715 26689
rect 10399 26624 10405 26688
rect 10469 26624 10485 26688
rect 10549 26624 10565 26688
rect 10629 26624 10645 26688
rect 10709 26624 10715 26688
rect 10399 26623 10715 26624
rect 16701 26688 17017 26689
rect 16701 26624 16707 26688
rect 16771 26624 16787 26688
rect 16851 26624 16867 26688
rect 16931 26624 16947 26688
rect 17011 26624 17017 26688
rect 16701 26623 17017 26624
rect 23003 26688 23319 26689
rect 23003 26624 23009 26688
rect 23073 26624 23089 26688
rect 23153 26624 23169 26688
rect 23233 26624 23249 26688
rect 23313 26624 23319 26688
rect 23003 26623 23319 26624
rect 4757 26144 5073 26145
rect 4757 26080 4763 26144
rect 4827 26080 4843 26144
rect 4907 26080 4923 26144
rect 4987 26080 5003 26144
rect 5067 26080 5073 26144
rect 4757 26079 5073 26080
rect 11059 26144 11375 26145
rect 11059 26080 11065 26144
rect 11129 26080 11145 26144
rect 11209 26080 11225 26144
rect 11289 26080 11305 26144
rect 11369 26080 11375 26144
rect 11059 26079 11375 26080
rect 17361 26144 17677 26145
rect 17361 26080 17367 26144
rect 17431 26080 17447 26144
rect 17511 26080 17527 26144
rect 17591 26080 17607 26144
rect 17671 26080 17677 26144
rect 17361 26079 17677 26080
rect 23663 26144 23979 26145
rect 23663 26080 23669 26144
rect 23733 26080 23749 26144
rect 23813 26080 23829 26144
rect 23893 26080 23909 26144
rect 23973 26080 23979 26144
rect 23663 26079 23979 26080
rect 4097 25600 4413 25601
rect 4097 25536 4103 25600
rect 4167 25536 4183 25600
rect 4247 25536 4263 25600
rect 4327 25536 4343 25600
rect 4407 25536 4413 25600
rect 4097 25535 4413 25536
rect 10399 25600 10715 25601
rect 10399 25536 10405 25600
rect 10469 25536 10485 25600
rect 10549 25536 10565 25600
rect 10629 25536 10645 25600
rect 10709 25536 10715 25600
rect 10399 25535 10715 25536
rect 16701 25600 17017 25601
rect 16701 25536 16707 25600
rect 16771 25536 16787 25600
rect 16851 25536 16867 25600
rect 16931 25536 16947 25600
rect 17011 25536 17017 25600
rect 16701 25535 17017 25536
rect 23003 25600 23319 25601
rect 23003 25536 23009 25600
rect 23073 25536 23089 25600
rect 23153 25536 23169 25600
rect 23233 25536 23249 25600
rect 23313 25536 23319 25600
rect 23003 25535 23319 25536
rect 0 25258 800 25288
rect 3233 25258 3299 25261
rect 0 25256 3299 25258
rect 0 25200 3238 25256
rect 3294 25200 3299 25256
rect 0 25198 3299 25200
rect 0 25168 800 25198
rect 3233 25195 3299 25198
rect 9121 25258 9187 25261
rect 10133 25258 10199 25261
rect 9121 25256 10199 25258
rect 9121 25200 9126 25256
rect 9182 25200 10138 25256
rect 10194 25200 10199 25256
rect 9121 25198 10199 25200
rect 9121 25195 9187 25198
rect 10133 25195 10199 25198
rect 25773 25258 25839 25261
rect 26681 25258 27481 25288
rect 25773 25256 27481 25258
rect 25773 25200 25778 25256
rect 25834 25200 27481 25256
rect 25773 25198 27481 25200
rect 25773 25195 25839 25198
rect 26681 25168 27481 25198
rect 4757 25056 5073 25057
rect 4757 24992 4763 25056
rect 4827 24992 4843 25056
rect 4907 24992 4923 25056
rect 4987 24992 5003 25056
rect 5067 24992 5073 25056
rect 4757 24991 5073 24992
rect 11059 25056 11375 25057
rect 11059 24992 11065 25056
rect 11129 24992 11145 25056
rect 11209 24992 11225 25056
rect 11289 24992 11305 25056
rect 11369 24992 11375 25056
rect 11059 24991 11375 24992
rect 17361 25056 17677 25057
rect 17361 24992 17367 25056
rect 17431 24992 17447 25056
rect 17511 24992 17527 25056
rect 17591 24992 17607 25056
rect 17671 24992 17677 25056
rect 17361 24991 17677 24992
rect 23663 25056 23979 25057
rect 23663 24992 23669 25056
rect 23733 24992 23749 25056
rect 23813 24992 23829 25056
rect 23893 24992 23909 25056
rect 23973 24992 23979 25056
rect 23663 24991 23979 24992
rect 17125 24850 17191 24853
rect 17769 24850 17835 24853
rect 17125 24848 17835 24850
rect 17125 24792 17130 24848
rect 17186 24792 17774 24848
rect 17830 24792 17835 24848
rect 17125 24790 17835 24792
rect 17125 24787 17191 24790
rect 17769 24787 17835 24790
rect 4097 24512 4413 24513
rect 4097 24448 4103 24512
rect 4167 24448 4183 24512
rect 4247 24448 4263 24512
rect 4327 24448 4343 24512
rect 4407 24448 4413 24512
rect 4097 24447 4413 24448
rect 10399 24512 10715 24513
rect 10399 24448 10405 24512
rect 10469 24448 10485 24512
rect 10549 24448 10565 24512
rect 10629 24448 10645 24512
rect 10709 24448 10715 24512
rect 10399 24447 10715 24448
rect 16701 24512 17017 24513
rect 16701 24448 16707 24512
rect 16771 24448 16787 24512
rect 16851 24448 16867 24512
rect 16931 24448 16947 24512
rect 17011 24448 17017 24512
rect 16701 24447 17017 24448
rect 23003 24512 23319 24513
rect 23003 24448 23009 24512
rect 23073 24448 23089 24512
rect 23153 24448 23169 24512
rect 23233 24448 23249 24512
rect 23313 24448 23319 24512
rect 23003 24447 23319 24448
rect 20253 24170 20319 24173
rect 23105 24170 23171 24173
rect 23749 24170 23815 24173
rect 20253 24168 23815 24170
rect 20253 24112 20258 24168
rect 20314 24112 23110 24168
rect 23166 24112 23754 24168
rect 23810 24112 23815 24168
rect 20253 24110 23815 24112
rect 20253 24107 20319 24110
rect 23105 24107 23171 24110
rect 23749 24107 23815 24110
rect 9949 24034 10015 24037
rect 10685 24034 10751 24037
rect 9949 24032 10751 24034
rect 9949 23976 9954 24032
rect 10010 23976 10690 24032
rect 10746 23976 10751 24032
rect 9949 23974 10751 23976
rect 9949 23971 10015 23974
rect 10685 23971 10751 23974
rect 4757 23968 5073 23969
rect 4757 23904 4763 23968
rect 4827 23904 4843 23968
rect 4907 23904 4923 23968
rect 4987 23904 5003 23968
rect 5067 23904 5073 23968
rect 4757 23903 5073 23904
rect 11059 23968 11375 23969
rect 11059 23904 11065 23968
rect 11129 23904 11145 23968
rect 11209 23904 11225 23968
rect 11289 23904 11305 23968
rect 11369 23904 11375 23968
rect 11059 23903 11375 23904
rect 17361 23968 17677 23969
rect 17361 23904 17367 23968
rect 17431 23904 17447 23968
rect 17511 23904 17527 23968
rect 17591 23904 17607 23968
rect 17671 23904 17677 23968
rect 17361 23903 17677 23904
rect 23663 23968 23979 23969
rect 23663 23904 23669 23968
rect 23733 23904 23749 23968
rect 23813 23904 23829 23968
rect 23893 23904 23909 23968
rect 23973 23904 23979 23968
rect 23663 23903 23979 23904
rect 9305 23898 9371 23901
rect 10041 23898 10107 23901
rect 9305 23896 10107 23898
rect 9305 23840 9310 23896
rect 9366 23840 10046 23896
rect 10102 23840 10107 23896
rect 9305 23838 10107 23840
rect 9305 23835 9371 23838
rect 10041 23835 10107 23838
rect 5165 23762 5231 23765
rect 27061 23762 27127 23765
rect 5165 23760 27127 23762
rect 5165 23704 5170 23760
rect 5226 23704 27066 23760
rect 27122 23704 27127 23760
rect 5165 23702 27127 23704
rect 5165 23699 5231 23702
rect 27061 23699 27127 23702
rect 6453 23626 6519 23629
rect 6821 23626 6887 23629
rect 11053 23626 11119 23629
rect 6453 23624 11119 23626
rect 6453 23568 6458 23624
rect 6514 23568 6826 23624
rect 6882 23568 11058 23624
rect 11114 23568 11119 23624
rect 6453 23566 11119 23568
rect 6453 23563 6519 23566
rect 6821 23563 6887 23566
rect 11053 23563 11119 23566
rect 5533 23492 5599 23493
rect 5533 23488 5580 23492
rect 5644 23490 5650 23492
rect 9489 23490 9555 23493
rect 10133 23490 10199 23493
rect 5533 23432 5538 23488
rect 5533 23428 5580 23432
rect 5644 23430 5690 23490
rect 9489 23488 10199 23490
rect 9489 23432 9494 23488
rect 9550 23432 10138 23488
rect 10194 23432 10199 23488
rect 9489 23430 10199 23432
rect 5644 23428 5650 23430
rect 5533 23427 5599 23428
rect 9489 23427 9555 23430
rect 10133 23427 10199 23430
rect 4097 23424 4413 23425
rect 4097 23360 4103 23424
rect 4167 23360 4183 23424
rect 4247 23360 4263 23424
rect 4327 23360 4343 23424
rect 4407 23360 4413 23424
rect 4097 23359 4413 23360
rect 10399 23424 10715 23425
rect 10399 23360 10405 23424
rect 10469 23360 10485 23424
rect 10549 23360 10565 23424
rect 10629 23360 10645 23424
rect 10709 23360 10715 23424
rect 10399 23359 10715 23360
rect 16701 23424 17017 23425
rect 16701 23360 16707 23424
rect 16771 23360 16787 23424
rect 16851 23360 16867 23424
rect 16931 23360 16947 23424
rect 17011 23360 17017 23424
rect 16701 23359 17017 23360
rect 23003 23424 23319 23425
rect 23003 23360 23009 23424
rect 23073 23360 23089 23424
rect 23153 23360 23169 23424
rect 23233 23360 23249 23424
rect 23313 23360 23319 23424
rect 23003 23359 23319 23360
rect 9949 23354 10015 23357
rect 20345 23354 20411 23357
rect 20713 23354 20779 23357
rect 9949 23352 10196 23354
rect 9949 23296 9954 23352
rect 10010 23296 10196 23352
rect 9949 23294 10196 23296
rect 9949 23291 10015 23294
rect 10136 23218 10196 23294
rect 20345 23352 20779 23354
rect 20345 23296 20350 23352
rect 20406 23296 20718 23352
rect 20774 23296 20779 23352
rect 20345 23294 20779 23296
rect 20345 23291 20411 23294
rect 20713 23291 20779 23294
rect 10777 23218 10843 23221
rect 10136 23216 10843 23218
rect 10136 23160 10782 23216
rect 10838 23160 10843 23216
rect 10136 23158 10843 23160
rect 10777 23155 10843 23158
rect 20069 23218 20135 23221
rect 20713 23218 20779 23221
rect 20069 23216 20779 23218
rect 20069 23160 20074 23216
rect 20130 23160 20718 23216
rect 20774 23160 20779 23216
rect 20069 23158 20779 23160
rect 20069 23155 20135 23158
rect 20713 23155 20779 23158
rect 19885 23082 19951 23085
rect 21265 23082 21331 23085
rect 19885 23080 21331 23082
rect 19885 23024 19890 23080
rect 19946 23024 21270 23080
rect 21326 23024 21331 23080
rect 19885 23022 21331 23024
rect 19885 23019 19951 23022
rect 21265 23019 21331 23022
rect 4757 22880 5073 22881
rect 4757 22816 4763 22880
rect 4827 22816 4843 22880
rect 4907 22816 4923 22880
rect 4987 22816 5003 22880
rect 5067 22816 5073 22880
rect 4757 22815 5073 22816
rect 11059 22880 11375 22881
rect 11059 22816 11065 22880
rect 11129 22816 11145 22880
rect 11209 22816 11225 22880
rect 11289 22816 11305 22880
rect 11369 22816 11375 22880
rect 11059 22815 11375 22816
rect 17361 22880 17677 22881
rect 17361 22816 17367 22880
rect 17431 22816 17447 22880
rect 17511 22816 17527 22880
rect 17591 22816 17607 22880
rect 17671 22816 17677 22880
rect 17361 22815 17677 22816
rect 23663 22880 23979 22881
rect 23663 22816 23669 22880
rect 23733 22816 23749 22880
rect 23813 22816 23829 22880
rect 23893 22816 23909 22880
rect 23973 22816 23979 22880
rect 23663 22815 23979 22816
rect 4097 22336 4413 22337
rect 4097 22272 4103 22336
rect 4167 22272 4183 22336
rect 4247 22272 4263 22336
rect 4327 22272 4343 22336
rect 4407 22272 4413 22336
rect 4097 22271 4413 22272
rect 10399 22336 10715 22337
rect 10399 22272 10405 22336
rect 10469 22272 10485 22336
rect 10549 22272 10565 22336
rect 10629 22272 10645 22336
rect 10709 22272 10715 22336
rect 10399 22271 10715 22272
rect 16701 22336 17017 22337
rect 16701 22272 16707 22336
rect 16771 22272 16787 22336
rect 16851 22272 16867 22336
rect 16931 22272 16947 22336
rect 17011 22272 17017 22336
rect 16701 22271 17017 22272
rect 23003 22336 23319 22337
rect 23003 22272 23009 22336
rect 23073 22272 23089 22336
rect 23153 22272 23169 22336
rect 23233 22272 23249 22336
rect 23313 22272 23319 22336
rect 23003 22271 23319 22272
rect 4153 21994 4219 21997
rect 4889 21994 4955 21997
rect 6126 21994 6132 21996
rect 4153 21992 6132 21994
rect 4153 21936 4158 21992
rect 4214 21936 4894 21992
rect 4950 21936 6132 21992
rect 4153 21934 6132 21936
rect 4153 21931 4219 21934
rect 4889 21931 4955 21934
rect 6126 21932 6132 21934
rect 6196 21932 6202 21996
rect 4757 21792 5073 21793
rect 4757 21728 4763 21792
rect 4827 21728 4843 21792
rect 4907 21728 4923 21792
rect 4987 21728 5003 21792
rect 5067 21728 5073 21792
rect 4757 21727 5073 21728
rect 11059 21792 11375 21793
rect 11059 21728 11065 21792
rect 11129 21728 11145 21792
rect 11209 21728 11225 21792
rect 11289 21728 11305 21792
rect 11369 21728 11375 21792
rect 11059 21727 11375 21728
rect 17361 21792 17677 21793
rect 17361 21728 17367 21792
rect 17431 21728 17447 21792
rect 17511 21728 17527 21792
rect 17591 21728 17607 21792
rect 17671 21728 17677 21792
rect 17361 21727 17677 21728
rect 23663 21792 23979 21793
rect 23663 21728 23669 21792
rect 23733 21728 23749 21792
rect 23813 21728 23829 21792
rect 23893 21728 23909 21792
rect 23973 21728 23979 21792
rect 23663 21727 23979 21728
rect 4097 21248 4413 21249
rect 0 21178 800 21208
rect 4097 21184 4103 21248
rect 4167 21184 4183 21248
rect 4247 21184 4263 21248
rect 4327 21184 4343 21248
rect 4407 21184 4413 21248
rect 4097 21183 4413 21184
rect 10399 21248 10715 21249
rect 10399 21184 10405 21248
rect 10469 21184 10485 21248
rect 10549 21184 10565 21248
rect 10629 21184 10645 21248
rect 10709 21184 10715 21248
rect 10399 21183 10715 21184
rect 16701 21248 17017 21249
rect 16701 21184 16707 21248
rect 16771 21184 16787 21248
rect 16851 21184 16867 21248
rect 16931 21184 16947 21248
rect 17011 21184 17017 21248
rect 16701 21183 17017 21184
rect 23003 21248 23319 21249
rect 23003 21184 23009 21248
rect 23073 21184 23089 21248
rect 23153 21184 23169 21248
rect 23233 21184 23249 21248
rect 23313 21184 23319 21248
rect 23003 21183 23319 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 25773 21178 25839 21181
rect 26681 21178 27481 21208
rect 25773 21176 27481 21178
rect 25773 21120 25778 21176
rect 25834 21120 27481 21176
rect 25773 21118 27481 21120
rect 25773 21115 25839 21118
rect 26681 21088 27481 21118
rect 14273 20906 14339 20909
rect 19057 20906 19123 20909
rect 19425 20906 19491 20909
rect 14273 20904 19491 20906
rect 14273 20848 14278 20904
rect 14334 20848 19062 20904
rect 19118 20848 19430 20904
rect 19486 20848 19491 20904
rect 14273 20846 19491 20848
rect 14273 20843 14339 20846
rect 19057 20843 19123 20846
rect 19425 20843 19491 20846
rect 4757 20704 5073 20705
rect 4757 20640 4763 20704
rect 4827 20640 4843 20704
rect 4907 20640 4923 20704
rect 4987 20640 5003 20704
rect 5067 20640 5073 20704
rect 4757 20639 5073 20640
rect 11059 20704 11375 20705
rect 11059 20640 11065 20704
rect 11129 20640 11145 20704
rect 11209 20640 11225 20704
rect 11289 20640 11305 20704
rect 11369 20640 11375 20704
rect 11059 20639 11375 20640
rect 17361 20704 17677 20705
rect 17361 20640 17367 20704
rect 17431 20640 17447 20704
rect 17511 20640 17527 20704
rect 17591 20640 17607 20704
rect 17671 20640 17677 20704
rect 17361 20639 17677 20640
rect 23663 20704 23979 20705
rect 23663 20640 23669 20704
rect 23733 20640 23749 20704
rect 23813 20640 23829 20704
rect 23893 20640 23909 20704
rect 23973 20640 23979 20704
rect 23663 20639 23979 20640
rect 1577 20498 1643 20501
rect 15193 20498 15259 20501
rect 1577 20496 15259 20498
rect 1577 20440 1582 20496
rect 1638 20440 15198 20496
rect 15254 20440 15259 20496
rect 1577 20438 15259 20440
rect 1577 20435 1643 20438
rect 15193 20435 15259 20438
rect 4097 20160 4413 20161
rect 4097 20096 4103 20160
rect 4167 20096 4183 20160
rect 4247 20096 4263 20160
rect 4327 20096 4343 20160
rect 4407 20096 4413 20160
rect 4097 20095 4413 20096
rect 10399 20160 10715 20161
rect 10399 20096 10405 20160
rect 10469 20096 10485 20160
rect 10549 20096 10565 20160
rect 10629 20096 10645 20160
rect 10709 20096 10715 20160
rect 10399 20095 10715 20096
rect 16701 20160 17017 20161
rect 16701 20096 16707 20160
rect 16771 20096 16787 20160
rect 16851 20096 16867 20160
rect 16931 20096 16947 20160
rect 17011 20096 17017 20160
rect 16701 20095 17017 20096
rect 23003 20160 23319 20161
rect 23003 20096 23009 20160
rect 23073 20096 23089 20160
rect 23153 20096 23169 20160
rect 23233 20096 23249 20160
rect 23313 20096 23319 20160
rect 23003 20095 23319 20096
rect 2589 19818 2655 19821
rect 17125 19818 17191 19821
rect 2589 19816 17191 19818
rect 2589 19760 2594 19816
rect 2650 19760 17130 19816
rect 17186 19760 17191 19816
rect 2589 19758 17191 19760
rect 2589 19755 2655 19758
rect 17125 19755 17191 19758
rect 4757 19616 5073 19617
rect 4757 19552 4763 19616
rect 4827 19552 4843 19616
rect 4907 19552 4923 19616
rect 4987 19552 5003 19616
rect 5067 19552 5073 19616
rect 4757 19551 5073 19552
rect 11059 19616 11375 19617
rect 11059 19552 11065 19616
rect 11129 19552 11145 19616
rect 11209 19552 11225 19616
rect 11289 19552 11305 19616
rect 11369 19552 11375 19616
rect 11059 19551 11375 19552
rect 17361 19616 17677 19617
rect 17361 19552 17367 19616
rect 17431 19552 17447 19616
rect 17511 19552 17527 19616
rect 17591 19552 17607 19616
rect 17671 19552 17677 19616
rect 17361 19551 17677 19552
rect 23663 19616 23979 19617
rect 23663 19552 23669 19616
rect 23733 19552 23749 19616
rect 23813 19552 23829 19616
rect 23893 19552 23909 19616
rect 23973 19552 23979 19616
rect 23663 19551 23979 19552
rect 4797 19410 4863 19413
rect 10317 19410 10383 19413
rect 4797 19408 10383 19410
rect 4797 19352 4802 19408
rect 4858 19352 10322 19408
rect 10378 19352 10383 19408
rect 4797 19350 10383 19352
rect 4797 19347 4863 19350
rect 10317 19347 10383 19350
rect 4097 19072 4413 19073
rect 4097 19008 4103 19072
rect 4167 19008 4183 19072
rect 4247 19008 4263 19072
rect 4327 19008 4343 19072
rect 4407 19008 4413 19072
rect 4097 19007 4413 19008
rect 10399 19072 10715 19073
rect 10399 19008 10405 19072
rect 10469 19008 10485 19072
rect 10549 19008 10565 19072
rect 10629 19008 10645 19072
rect 10709 19008 10715 19072
rect 10399 19007 10715 19008
rect 16701 19072 17017 19073
rect 16701 19008 16707 19072
rect 16771 19008 16787 19072
rect 16851 19008 16867 19072
rect 16931 19008 16947 19072
rect 17011 19008 17017 19072
rect 16701 19007 17017 19008
rect 23003 19072 23319 19073
rect 23003 19008 23009 19072
rect 23073 19008 23089 19072
rect 23153 19008 23169 19072
rect 23233 19008 23249 19072
rect 23313 19008 23319 19072
rect 23003 19007 23319 19008
rect 14457 18866 14523 18869
rect 22737 18866 22803 18869
rect 14457 18864 22803 18866
rect 14457 18808 14462 18864
rect 14518 18808 22742 18864
rect 22798 18808 22803 18864
rect 14457 18806 22803 18808
rect 14457 18803 14523 18806
rect 22737 18803 22803 18806
rect 4757 18528 5073 18529
rect 4757 18464 4763 18528
rect 4827 18464 4843 18528
rect 4907 18464 4923 18528
rect 4987 18464 5003 18528
rect 5067 18464 5073 18528
rect 4757 18463 5073 18464
rect 11059 18528 11375 18529
rect 11059 18464 11065 18528
rect 11129 18464 11145 18528
rect 11209 18464 11225 18528
rect 11289 18464 11305 18528
rect 11369 18464 11375 18528
rect 11059 18463 11375 18464
rect 17361 18528 17677 18529
rect 17361 18464 17367 18528
rect 17431 18464 17447 18528
rect 17511 18464 17527 18528
rect 17591 18464 17607 18528
rect 17671 18464 17677 18528
rect 17361 18463 17677 18464
rect 23663 18528 23979 18529
rect 23663 18464 23669 18528
rect 23733 18464 23749 18528
rect 23813 18464 23829 18528
rect 23893 18464 23909 18528
rect 23973 18464 23979 18528
rect 23663 18463 23979 18464
rect 16389 18458 16455 18461
rect 17217 18458 17283 18461
rect 16389 18456 17283 18458
rect 16389 18400 16394 18456
rect 16450 18400 17222 18456
rect 17278 18400 17283 18456
rect 16389 18398 17283 18400
rect 16389 18395 16455 18398
rect 17217 18395 17283 18398
rect 14641 18322 14707 18325
rect 25221 18322 25287 18325
rect 14641 18320 25287 18322
rect 14641 18264 14646 18320
rect 14702 18264 25226 18320
rect 25282 18264 25287 18320
rect 14641 18262 25287 18264
rect 14641 18259 14707 18262
rect 25221 18259 25287 18262
rect 16113 18186 16179 18189
rect 17401 18186 17467 18189
rect 16113 18184 17467 18186
rect 16113 18128 16118 18184
rect 16174 18128 17406 18184
rect 17462 18128 17467 18184
rect 16113 18126 17467 18128
rect 16113 18123 16179 18126
rect 17401 18123 17467 18126
rect 4097 17984 4413 17985
rect 4097 17920 4103 17984
rect 4167 17920 4183 17984
rect 4247 17920 4263 17984
rect 4327 17920 4343 17984
rect 4407 17920 4413 17984
rect 4097 17919 4413 17920
rect 10399 17984 10715 17985
rect 10399 17920 10405 17984
rect 10469 17920 10485 17984
rect 10549 17920 10565 17984
rect 10629 17920 10645 17984
rect 10709 17920 10715 17984
rect 10399 17919 10715 17920
rect 16701 17984 17017 17985
rect 16701 17920 16707 17984
rect 16771 17920 16787 17984
rect 16851 17920 16867 17984
rect 16931 17920 16947 17984
rect 17011 17920 17017 17984
rect 16701 17919 17017 17920
rect 23003 17984 23319 17985
rect 23003 17920 23009 17984
rect 23073 17920 23089 17984
rect 23153 17920 23169 17984
rect 23233 17920 23249 17984
rect 23313 17920 23319 17984
rect 23003 17919 23319 17920
rect 7925 17914 7991 17917
rect 10133 17914 10199 17917
rect 7925 17912 10199 17914
rect 7925 17856 7930 17912
rect 7986 17856 10138 17912
rect 10194 17856 10199 17912
rect 7925 17854 10199 17856
rect 7925 17851 7991 17854
rect 10133 17851 10199 17854
rect 6126 17444 6132 17508
rect 6196 17506 6202 17508
rect 6637 17506 6703 17509
rect 6196 17504 6703 17506
rect 6196 17448 6642 17504
rect 6698 17448 6703 17504
rect 6196 17446 6703 17448
rect 6196 17444 6202 17446
rect 6637 17443 6703 17446
rect 4757 17440 5073 17441
rect 4757 17376 4763 17440
rect 4827 17376 4843 17440
rect 4907 17376 4923 17440
rect 4987 17376 5003 17440
rect 5067 17376 5073 17440
rect 4757 17375 5073 17376
rect 11059 17440 11375 17441
rect 11059 17376 11065 17440
rect 11129 17376 11145 17440
rect 11209 17376 11225 17440
rect 11289 17376 11305 17440
rect 11369 17376 11375 17440
rect 11059 17375 11375 17376
rect 17361 17440 17677 17441
rect 17361 17376 17367 17440
rect 17431 17376 17447 17440
rect 17511 17376 17527 17440
rect 17591 17376 17607 17440
rect 17671 17376 17677 17440
rect 17361 17375 17677 17376
rect 23663 17440 23979 17441
rect 23663 17376 23669 17440
rect 23733 17376 23749 17440
rect 23813 17376 23829 17440
rect 23893 17376 23909 17440
rect 23973 17376 23979 17440
rect 23663 17375 23979 17376
rect 25865 17098 25931 17101
rect 26681 17098 27481 17128
rect 25865 17096 27481 17098
rect 25865 17040 25870 17096
rect 25926 17040 27481 17096
rect 25865 17038 27481 17040
rect 25865 17035 25931 17038
rect 26681 17008 27481 17038
rect 4097 16896 4413 16897
rect 4097 16832 4103 16896
rect 4167 16832 4183 16896
rect 4247 16832 4263 16896
rect 4327 16832 4343 16896
rect 4407 16832 4413 16896
rect 4097 16831 4413 16832
rect 10399 16896 10715 16897
rect 10399 16832 10405 16896
rect 10469 16832 10485 16896
rect 10549 16832 10565 16896
rect 10629 16832 10645 16896
rect 10709 16832 10715 16896
rect 10399 16831 10715 16832
rect 16701 16896 17017 16897
rect 16701 16832 16707 16896
rect 16771 16832 16787 16896
rect 16851 16832 16867 16896
rect 16931 16832 16947 16896
rect 17011 16832 17017 16896
rect 16701 16831 17017 16832
rect 23003 16896 23319 16897
rect 23003 16832 23009 16896
rect 23073 16832 23089 16896
rect 23153 16832 23169 16896
rect 23233 16832 23249 16896
rect 23313 16832 23319 16896
rect 23003 16831 23319 16832
rect 20253 16690 20319 16693
rect 23197 16690 23263 16693
rect 20253 16688 23263 16690
rect 20253 16632 20258 16688
rect 20314 16632 23202 16688
rect 23258 16632 23263 16688
rect 20253 16630 23263 16632
rect 20253 16627 20319 16630
rect 23197 16627 23263 16630
rect 20713 16554 20779 16557
rect 21265 16554 21331 16557
rect 20713 16552 21331 16554
rect 20713 16496 20718 16552
rect 20774 16496 21270 16552
rect 21326 16496 21331 16552
rect 20713 16494 21331 16496
rect 20713 16491 20779 16494
rect 21265 16491 21331 16494
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 4757 16352 5073 16353
rect 4757 16288 4763 16352
rect 4827 16288 4843 16352
rect 4907 16288 4923 16352
rect 4987 16288 5003 16352
rect 5067 16288 5073 16352
rect 4757 16287 5073 16288
rect 11059 16352 11375 16353
rect 11059 16288 11065 16352
rect 11129 16288 11145 16352
rect 11209 16288 11225 16352
rect 11289 16288 11305 16352
rect 11369 16288 11375 16352
rect 11059 16287 11375 16288
rect 17361 16352 17677 16353
rect 17361 16288 17367 16352
rect 17431 16288 17447 16352
rect 17511 16288 17527 16352
rect 17591 16288 17607 16352
rect 17671 16288 17677 16352
rect 17361 16287 17677 16288
rect 23663 16352 23979 16353
rect 23663 16288 23669 16352
rect 23733 16288 23749 16352
rect 23813 16288 23829 16352
rect 23893 16288 23909 16352
rect 23973 16288 23979 16352
rect 23663 16287 23979 16288
rect 4097 15808 4413 15809
rect 4097 15744 4103 15808
rect 4167 15744 4183 15808
rect 4247 15744 4263 15808
rect 4327 15744 4343 15808
rect 4407 15744 4413 15808
rect 4097 15743 4413 15744
rect 10399 15808 10715 15809
rect 10399 15744 10405 15808
rect 10469 15744 10485 15808
rect 10549 15744 10565 15808
rect 10629 15744 10645 15808
rect 10709 15744 10715 15808
rect 10399 15743 10715 15744
rect 16701 15808 17017 15809
rect 16701 15744 16707 15808
rect 16771 15744 16787 15808
rect 16851 15744 16867 15808
rect 16931 15744 16947 15808
rect 17011 15744 17017 15808
rect 16701 15743 17017 15744
rect 23003 15808 23319 15809
rect 23003 15744 23009 15808
rect 23073 15744 23089 15808
rect 23153 15744 23169 15808
rect 23233 15744 23249 15808
rect 23313 15744 23319 15808
rect 23003 15743 23319 15744
rect 4757 15264 5073 15265
rect 4757 15200 4763 15264
rect 4827 15200 4843 15264
rect 4907 15200 4923 15264
rect 4987 15200 5003 15264
rect 5067 15200 5073 15264
rect 4757 15199 5073 15200
rect 11059 15264 11375 15265
rect 11059 15200 11065 15264
rect 11129 15200 11145 15264
rect 11209 15200 11225 15264
rect 11289 15200 11305 15264
rect 11369 15200 11375 15264
rect 11059 15199 11375 15200
rect 17361 15264 17677 15265
rect 17361 15200 17367 15264
rect 17431 15200 17447 15264
rect 17511 15200 17527 15264
rect 17591 15200 17607 15264
rect 17671 15200 17677 15264
rect 17361 15199 17677 15200
rect 23663 15264 23979 15265
rect 23663 15200 23669 15264
rect 23733 15200 23749 15264
rect 23813 15200 23829 15264
rect 23893 15200 23909 15264
rect 23973 15200 23979 15264
rect 23663 15199 23979 15200
rect 5574 14996 5580 15060
rect 5644 15058 5650 15060
rect 12617 15058 12683 15061
rect 5644 15056 12683 15058
rect 5644 15000 12622 15056
rect 12678 15000 12683 15056
rect 5644 14998 12683 15000
rect 5644 14996 5650 14998
rect 12617 14995 12683 14998
rect 4097 14720 4413 14721
rect 4097 14656 4103 14720
rect 4167 14656 4183 14720
rect 4247 14656 4263 14720
rect 4327 14656 4343 14720
rect 4407 14656 4413 14720
rect 4097 14655 4413 14656
rect 10399 14720 10715 14721
rect 10399 14656 10405 14720
rect 10469 14656 10485 14720
rect 10549 14656 10565 14720
rect 10629 14656 10645 14720
rect 10709 14656 10715 14720
rect 10399 14655 10715 14656
rect 16701 14720 17017 14721
rect 16701 14656 16707 14720
rect 16771 14656 16787 14720
rect 16851 14656 16867 14720
rect 16931 14656 16947 14720
rect 17011 14656 17017 14720
rect 16701 14655 17017 14656
rect 23003 14720 23319 14721
rect 23003 14656 23009 14720
rect 23073 14656 23089 14720
rect 23153 14656 23169 14720
rect 23233 14656 23249 14720
rect 23313 14656 23319 14720
rect 23003 14655 23319 14656
rect 4757 14176 5073 14177
rect 4757 14112 4763 14176
rect 4827 14112 4843 14176
rect 4907 14112 4923 14176
rect 4987 14112 5003 14176
rect 5067 14112 5073 14176
rect 4757 14111 5073 14112
rect 11059 14176 11375 14177
rect 11059 14112 11065 14176
rect 11129 14112 11145 14176
rect 11209 14112 11225 14176
rect 11289 14112 11305 14176
rect 11369 14112 11375 14176
rect 11059 14111 11375 14112
rect 17361 14176 17677 14177
rect 17361 14112 17367 14176
rect 17431 14112 17447 14176
rect 17511 14112 17527 14176
rect 17591 14112 17607 14176
rect 17671 14112 17677 14176
rect 17361 14111 17677 14112
rect 23663 14176 23979 14177
rect 23663 14112 23669 14176
rect 23733 14112 23749 14176
rect 23813 14112 23829 14176
rect 23893 14112 23909 14176
rect 23973 14112 23979 14176
rect 23663 14111 23979 14112
rect 4097 13632 4413 13633
rect 4097 13568 4103 13632
rect 4167 13568 4183 13632
rect 4247 13568 4263 13632
rect 4327 13568 4343 13632
rect 4407 13568 4413 13632
rect 4097 13567 4413 13568
rect 10399 13632 10715 13633
rect 10399 13568 10405 13632
rect 10469 13568 10485 13632
rect 10549 13568 10565 13632
rect 10629 13568 10645 13632
rect 10709 13568 10715 13632
rect 10399 13567 10715 13568
rect 16701 13632 17017 13633
rect 16701 13568 16707 13632
rect 16771 13568 16787 13632
rect 16851 13568 16867 13632
rect 16931 13568 16947 13632
rect 17011 13568 17017 13632
rect 16701 13567 17017 13568
rect 23003 13632 23319 13633
rect 23003 13568 23009 13632
rect 23073 13568 23089 13632
rect 23153 13568 23169 13632
rect 23233 13568 23249 13632
rect 23313 13568 23319 13632
rect 23003 13567 23319 13568
rect 4757 13088 5073 13089
rect 4757 13024 4763 13088
rect 4827 13024 4843 13088
rect 4907 13024 4923 13088
rect 4987 13024 5003 13088
rect 5067 13024 5073 13088
rect 4757 13023 5073 13024
rect 11059 13088 11375 13089
rect 11059 13024 11065 13088
rect 11129 13024 11145 13088
rect 11209 13024 11225 13088
rect 11289 13024 11305 13088
rect 11369 13024 11375 13088
rect 11059 13023 11375 13024
rect 17361 13088 17677 13089
rect 17361 13024 17367 13088
rect 17431 13024 17447 13088
rect 17511 13024 17527 13088
rect 17591 13024 17607 13088
rect 17671 13024 17677 13088
rect 17361 13023 17677 13024
rect 23663 13088 23979 13089
rect 23663 13024 23669 13088
rect 23733 13024 23749 13088
rect 23813 13024 23829 13088
rect 23893 13024 23909 13088
rect 23973 13024 23979 13088
rect 23663 13023 23979 13024
rect 25773 13018 25839 13021
rect 26681 13018 27481 13048
rect 25773 13016 27481 13018
rect 25773 12960 25778 13016
rect 25834 12960 27481 13016
rect 25773 12958 27481 12960
rect 25773 12955 25839 12958
rect 26681 12928 27481 12958
rect 4097 12544 4413 12545
rect 4097 12480 4103 12544
rect 4167 12480 4183 12544
rect 4247 12480 4263 12544
rect 4327 12480 4343 12544
rect 4407 12480 4413 12544
rect 4097 12479 4413 12480
rect 10399 12544 10715 12545
rect 10399 12480 10405 12544
rect 10469 12480 10485 12544
rect 10549 12480 10565 12544
rect 10629 12480 10645 12544
rect 10709 12480 10715 12544
rect 10399 12479 10715 12480
rect 16701 12544 17017 12545
rect 16701 12480 16707 12544
rect 16771 12480 16787 12544
rect 16851 12480 16867 12544
rect 16931 12480 16947 12544
rect 17011 12480 17017 12544
rect 16701 12479 17017 12480
rect 23003 12544 23319 12545
rect 23003 12480 23009 12544
rect 23073 12480 23089 12544
rect 23153 12480 23169 12544
rect 23233 12480 23249 12544
rect 23313 12480 23319 12544
rect 23003 12479 23319 12480
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 5441 12338 5507 12341
rect 5625 12338 5691 12341
rect 5441 12336 5691 12338
rect 5441 12280 5446 12336
rect 5502 12280 5630 12336
rect 5686 12280 5691 12336
rect 5441 12278 5691 12280
rect 5441 12275 5507 12278
rect 5625 12275 5691 12278
rect 4337 12202 4403 12205
rect 6821 12202 6887 12205
rect 8201 12202 8267 12205
rect 4337 12200 8267 12202
rect 4337 12144 4342 12200
rect 4398 12144 6826 12200
rect 6882 12144 8206 12200
rect 8262 12144 8267 12200
rect 4337 12142 8267 12144
rect 4337 12139 4403 12142
rect 6821 12139 6887 12142
rect 8201 12139 8267 12142
rect 4757 12000 5073 12001
rect 4757 11936 4763 12000
rect 4827 11936 4843 12000
rect 4907 11936 4923 12000
rect 4987 11936 5003 12000
rect 5067 11936 5073 12000
rect 4757 11935 5073 11936
rect 11059 12000 11375 12001
rect 11059 11936 11065 12000
rect 11129 11936 11145 12000
rect 11209 11936 11225 12000
rect 11289 11936 11305 12000
rect 11369 11936 11375 12000
rect 11059 11935 11375 11936
rect 17361 12000 17677 12001
rect 17361 11936 17367 12000
rect 17431 11936 17447 12000
rect 17511 11936 17527 12000
rect 17591 11936 17607 12000
rect 17671 11936 17677 12000
rect 17361 11935 17677 11936
rect 23663 12000 23979 12001
rect 23663 11936 23669 12000
rect 23733 11936 23749 12000
rect 23813 11936 23829 12000
rect 23893 11936 23909 12000
rect 23973 11936 23979 12000
rect 23663 11935 23979 11936
rect 4705 11794 4771 11797
rect 5349 11794 5415 11797
rect 4705 11792 5415 11794
rect 4705 11736 4710 11792
rect 4766 11736 5354 11792
rect 5410 11736 5415 11792
rect 4705 11734 5415 11736
rect 4705 11731 4771 11734
rect 5349 11731 5415 11734
rect 5533 11794 5599 11797
rect 6729 11794 6795 11797
rect 5533 11792 6795 11794
rect 5533 11736 5538 11792
rect 5594 11736 6734 11792
rect 6790 11736 6795 11792
rect 5533 11734 6795 11736
rect 5533 11731 5599 11734
rect 6729 11731 6795 11734
rect 20713 11794 20779 11797
rect 23105 11794 23171 11797
rect 20713 11792 23171 11794
rect 20713 11736 20718 11792
rect 20774 11736 23110 11792
rect 23166 11736 23171 11792
rect 20713 11734 23171 11736
rect 20713 11731 20779 11734
rect 23105 11731 23171 11734
rect 5625 11658 5691 11661
rect 6729 11658 6795 11661
rect 5625 11656 6795 11658
rect 5625 11600 5630 11656
rect 5686 11600 6734 11656
rect 6790 11600 6795 11656
rect 5625 11598 6795 11600
rect 5625 11595 5691 11598
rect 6729 11595 6795 11598
rect 4097 11456 4413 11457
rect 4097 11392 4103 11456
rect 4167 11392 4183 11456
rect 4247 11392 4263 11456
rect 4327 11392 4343 11456
rect 4407 11392 4413 11456
rect 4097 11391 4413 11392
rect 10399 11456 10715 11457
rect 10399 11392 10405 11456
rect 10469 11392 10485 11456
rect 10549 11392 10565 11456
rect 10629 11392 10645 11456
rect 10709 11392 10715 11456
rect 10399 11391 10715 11392
rect 16701 11456 17017 11457
rect 16701 11392 16707 11456
rect 16771 11392 16787 11456
rect 16851 11392 16867 11456
rect 16931 11392 16947 11456
rect 17011 11392 17017 11456
rect 16701 11391 17017 11392
rect 23003 11456 23319 11457
rect 23003 11392 23009 11456
rect 23073 11392 23089 11456
rect 23153 11392 23169 11456
rect 23233 11392 23249 11456
rect 23313 11392 23319 11456
rect 23003 11391 23319 11392
rect 5533 11252 5599 11253
rect 6361 11252 6427 11253
rect 5533 11248 5580 11252
rect 5644 11250 5650 11252
rect 5533 11192 5538 11248
rect 5533 11188 5580 11192
rect 5644 11190 5690 11250
rect 5644 11188 5650 11190
rect 6310 11188 6316 11252
rect 6380 11250 6427 11252
rect 6380 11248 6472 11250
rect 6422 11192 6472 11248
rect 6380 11190 6472 11192
rect 6380 11188 6427 11190
rect 5533 11187 5599 11188
rect 6361 11187 6427 11188
rect 6269 11114 6335 11117
rect 7649 11114 7715 11117
rect 6269 11112 7715 11114
rect 6269 11056 6274 11112
rect 6330 11056 7654 11112
rect 7710 11056 7715 11112
rect 6269 11054 7715 11056
rect 6269 11051 6335 11054
rect 7649 11051 7715 11054
rect 4757 10912 5073 10913
rect 4757 10848 4763 10912
rect 4827 10848 4843 10912
rect 4907 10848 4923 10912
rect 4987 10848 5003 10912
rect 5067 10848 5073 10912
rect 4757 10847 5073 10848
rect 11059 10912 11375 10913
rect 11059 10848 11065 10912
rect 11129 10848 11145 10912
rect 11209 10848 11225 10912
rect 11289 10848 11305 10912
rect 11369 10848 11375 10912
rect 11059 10847 11375 10848
rect 17361 10912 17677 10913
rect 17361 10848 17367 10912
rect 17431 10848 17447 10912
rect 17511 10848 17527 10912
rect 17591 10848 17607 10912
rect 17671 10848 17677 10912
rect 17361 10847 17677 10848
rect 23663 10912 23979 10913
rect 23663 10848 23669 10912
rect 23733 10848 23749 10912
rect 23813 10848 23829 10912
rect 23893 10848 23909 10912
rect 23973 10848 23979 10912
rect 23663 10847 23979 10848
rect 4097 10368 4413 10369
rect 4097 10304 4103 10368
rect 4167 10304 4183 10368
rect 4247 10304 4263 10368
rect 4327 10304 4343 10368
rect 4407 10304 4413 10368
rect 4097 10303 4413 10304
rect 10399 10368 10715 10369
rect 10399 10304 10405 10368
rect 10469 10304 10485 10368
rect 10549 10304 10565 10368
rect 10629 10304 10645 10368
rect 10709 10304 10715 10368
rect 10399 10303 10715 10304
rect 16701 10368 17017 10369
rect 16701 10304 16707 10368
rect 16771 10304 16787 10368
rect 16851 10304 16867 10368
rect 16931 10304 16947 10368
rect 17011 10304 17017 10368
rect 16701 10303 17017 10304
rect 23003 10368 23319 10369
rect 23003 10304 23009 10368
rect 23073 10304 23089 10368
rect 23153 10304 23169 10368
rect 23233 10304 23249 10368
rect 23313 10304 23319 10368
rect 23003 10303 23319 10304
rect 4757 9824 5073 9825
rect 4757 9760 4763 9824
rect 4827 9760 4843 9824
rect 4907 9760 4923 9824
rect 4987 9760 5003 9824
rect 5067 9760 5073 9824
rect 4757 9759 5073 9760
rect 11059 9824 11375 9825
rect 11059 9760 11065 9824
rect 11129 9760 11145 9824
rect 11209 9760 11225 9824
rect 11289 9760 11305 9824
rect 11369 9760 11375 9824
rect 11059 9759 11375 9760
rect 17361 9824 17677 9825
rect 17361 9760 17367 9824
rect 17431 9760 17447 9824
rect 17511 9760 17527 9824
rect 17591 9760 17607 9824
rect 17671 9760 17677 9824
rect 17361 9759 17677 9760
rect 23663 9824 23979 9825
rect 23663 9760 23669 9824
rect 23733 9760 23749 9824
rect 23813 9760 23829 9824
rect 23893 9760 23909 9824
rect 23973 9760 23979 9824
rect 23663 9759 23979 9760
rect 4097 9280 4413 9281
rect 4097 9216 4103 9280
rect 4167 9216 4183 9280
rect 4247 9216 4263 9280
rect 4327 9216 4343 9280
rect 4407 9216 4413 9280
rect 4097 9215 4413 9216
rect 10399 9280 10715 9281
rect 10399 9216 10405 9280
rect 10469 9216 10485 9280
rect 10549 9216 10565 9280
rect 10629 9216 10645 9280
rect 10709 9216 10715 9280
rect 10399 9215 10715 9216
rect 16701 9280 17017 9281
rect 16701 9216 16707 9280
rect 16771 9216 16787 9280
rect 16851 9216 16867 9280
rect 16931 9216 16947 9280
rect 17011 9216 17017 9280
rect 16701 9215 17017 9216
rect 23003 9280 23319 9281
rect 23003 9216 23009 9280
rect 23073 9216 23089 9280
rect 23153 9216 23169 9280
rect 23233 9216 23249 9280
rect 23313 9216 23319 9280
rect 23003 9215 23319 9216
rect 4797 9074 4863 9077
rect 6453 9074 6519 9077
rect 4797 9072 6519 9074
rect 4797 9016 4802 9072
rect 4858 9016 6458 9072
rect 6514 9016 6519 9072
rect 4797 9014 6519 9016
rect 4797 9011 4863 9014
rect 6453 9011 6519 9014
rect 15101 9074 15167 9077
rect 18781 9074 18847 9077
rect 15101 9072 18847 9074
rect 15101 9016 15106 9072
rect 15162 9016 18786 9072
rect 18842 9016 18847 9072
rect 15101 9014 18847 9016
rect 15101 9011 15167 9014
rect 18781 9011 18847 9014
rect 4889 8938 4955 8941
rect 4889 8936 5274 8938
rect 4889 8880 4894 8936
rect 4950 8880 5274 8936
rect 4889 8878 5274 8880
rect 4889 8875 4955 8878
rect 4757 8736 5073 8737
rect 4757 8672 4763 8736
rect 4827 8672 4843 8736
rect 4907 8672 4923 8736
rect 4987 8672 5003 8736
rect 5067 8672 5073 8736
rect 4757 8671 5073 8672
rect 4981 8530 5047 8533
rect 5214 8530 5274 8878
rect 11059 8736 11375 8737
rect 11059 8672 11065 8736
rect 11129 8672 11145 8736
rect 11209 8672 11225 8736
rect 11289 8672 11305 8736
rect 11369 8672 11375 8736
rect 11059 8671 11375 8672
rect 17361 8736 17677 8737
rect 17361 8672 17367 8736
rect 17431 8672 17447 8736
rect 17511 8672 17527 8736
rect 17591 8672 17607 8736
rect 17671 8672 17677 8736
rect 17361 8671 17677 8672
rect 23663 8736 23979 8737
rect 23663 8672 23669 8736
rect 23733 8672 23749 8736
rect 23813 8672 23829 8736
rect 23893 8672 23909 8736
rect 23973 8672 23979 8736
rect 23663 8671 23979 8672
rect 5533 8666 5599 8669
rect 6310 8666 6316 8668
rect 5533 8664 6316 8666
rect 5533 8608 5538 8664
rect 5594 8608 6316 8664
rect 5533 8606 6316 8608
rect 5533 8603 5599 8606
rect 6310 8604 6316 8606
rect 6380 8604 6386 8668
rect 4981 8528 5274 8530
rect 4981 8472 4986 8528
rect 5042 8472 5274 8528
rect 4981 8470 5274 8472
rect 4981 8467 5047 8470
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 25865 8258 25931 8261
rect 26681 8258 27481 8288
rect 25865 8256 27481 8258
rect 25865 8200 25870 8256
rect 25926 8200 27481 8256
rect 25865 8198 27481 8200
rect 25865 8195 25931 8198
rect 4097 8192 4413 8193
rect 4097 8128 4103 8192
rect 4167 8128 4183 8192
rect 4247 8128 4263 8192
rect 4327 8128 4343 8192
rect 4407 8128 4413 8192
rect 4097 8127 4413 8128
rect 10399 8192 10715 8193
rect 10399 8128 10405 8192
rect 10469 8128 10485 8192
rect 10549 8128 10565 8192
rect 10629 8128 10645 8192
rect 10709 8128 10715 8192
rect 10399 8127 10715 8128
rect 16701 8192 17017 8193
rect 16701 8128 16707 8192
rect 16771 8128 16787 8192
rect 16851 8128 16867 8192
rect 16931 8128 16947 8192
rect 17011 8128 17017 8192
rect 16701 8127 17017 8128
rect 23003 8192 23319 8193
rect 23003 8128 23009 8192
rect 23073 8128 23089 8192
rect 23153 8128 23169 8192
rect 23233 8128 23249 8192
rect 23313 8128 23319 8192
rect 26681 8168 27481 8198
rect 23003 8127 23319 8128
rect 5625 8124 5691 8125
rect 5574 8060 5580 8124
rect 5644 8122 5691 8124
rect 5644 8120 5736 8122
rect 5686 8064 5736 8120
rect 5644 8062 5736 8064
rect 5644 8060 5691 8062
rect 5625 8059 5691 8060
rect 4757 7648 5073 7649
rect 4757 7584 4763 7648
rect 4827 7584 4843 7648
rect 4907 7584 4923 7648
rect 4987 7584 5003 7648
rect 5067 7584 5073 7648
rect 4757 7583 5073 7584
rect 11059 7648 11375 7649
rect 11059 7584 11065 7648
rect 11129 7584 11145 7648
rect 11209 7584 11225 7648
rect 11289 7584 11305 7648
rect 11369 7584 11375 7648
rect 11059 7583 11375 7584
rect 17361 7648 17677 7649
rect 17361 7584 17367 7648
rect 17431 7584 17447 7648
rect 17511 7584 17527 7648
rect 17591 7584 17607 7648
rect 17671 7584 17677 7648
rect 17361 7583 17677 7584
rect 23663 7648 23979 7649
rect 23663 7584 23669 7648
rect 23733 7584 23749 7648
rect 23813 7584 23829 7648
rect 23893 7584 23909 7648
rect 23973 7584 23979 7648
rect 23663 7583 23979 7584
rect 4097 7104 4413 7105
rect 4097 7040 4103 7104
rect 4167 7040 4183 7104
rect 4247 7040 4263 7104
rect 4327 7040 4343 7104
rect 4407 7040 4413 7104
rect 4097 7039 4413 7040
rect 10399 7104 10715 7105
rect 10399 7040 10405 7104
rect 10469 7040 10485 7104
rect 10549 7040 10565 7104
rect 10629 7040 10645 7104
rect 10709 7040 10715 7104
rect 10399 7039 10715 7040
rect 16701 7104 17017 7105
rect 16701 7040 16707 7104
rect 16771 7040 16787 7104
rect 16851 7040 16867 7104
rect 16931 7040 16947 7104
rect 17011 7040 17017 7104
rect 16701 7039 17017 7040
rect 23003 7104 23319 7105
rect 23003 7040 23009 7104
rect 23073 7040 23089 7104
rect 23153 7040 23169 7104
rect 23233 7040 23249 7104
rect 23313 7040 23319 7104
rect 23003 7039 23319 7040
rect 4757 6560 5073 6561
rect 4757 6496 4763 6560
rect 4827 6496 4843 6560
rect 4907 6496 4923 6560
rect 4987 6496 5003 6560
rect 5067 6496 5073 6560
rect 4757 6495 5073 6496
rect 11059 6560 11375 6561
rect 11059 6496 11065 6560
rect 11129 6496 11145 6560
rect 11209 6496 11225 6560
rect 11289 6496 11305 6560
rect 11369 6496 11375 6560
rect 11059 6495 11375 6496
rect 17361 6560 17677 6561
rect 17361 6496 17367 6560
rect 17431 6496 17447 6560
rect 17511 6496 17527 6560
rect 17591 6496 17607 6560
rect 17671 6496 17677 6560
rect 17361 6495 17677 6496
rect 23663 6560 23979 6561
rect 23663 6496 23669 6560
rect 23733 6496 23749 6560
rect 23813 6496 23829 6560
rect 23893 6496 23909 6560
rect 23973 6496 23979 6560
rect 23663 6495 23979 6496
rect 19701 6354 19767 6357
rect 20805 6354 20871 6357
rect 19701 6352 20871 6354
rect 19701 6296 19706 6352
rect 19762 6296 20810 6352
rect 20866 6296 20871 6352
rect 19701 6294 20871 6296
rect 19701 6291 19767 6294
rect 20805 6291 20871 6294
rect 19333 6218 19399 6221
rect 20345 6218 20411 6221
rect 19333 6216 20411 6218
rect 19333 6160 19338 6216
rect 19394 6160 20350 6216
rect 20406 6160 20411 6216
rect 19333 6158 20411 6160
rect 19333 6155 19399 6158
rect 20345 6155 20411 6158
rect 19701 6082 19767 6085
rect 20529 6082 20595 6085
rect 22369 6082 22435 6085
rect 19701 6080 22435 6082
rect 19701 6024 19706 6080
rect 19762 6024 20534 6080
rect 20590 6024 22374 6080
rect 22430 6024 22435 6080
rect 19701 6022 22435 6024
rect 19701 6019 19767 6022
rect 20529 6019 20595 6022
rect 22369 6019 22435 6022
rect 4097 6016 4413 6017
rect 4097 5952 4103 6016
rect 4167 5952 4183 6016
rect 4247 5952 4263 6016
rect 4327 5952 4343 6016
rect 4407 5952 4413 6016
rect 4097 5951 4413 5952
rect 10399 6016 10715 6017
rect 10399 5952 10405 6016
rect 10469 5952 10485 6016
rect 10549 5952 10565 6016
rect 10629 5952 10645 6016
rect 10709 5952 10715 6016
rect 10399 5951 10715 5952
rect 16701 6016 17017 6017
rect 16701 5952 16707 6016
rect 16771 5952 16787 6016
rect 16851 5952 16867 6016
rect 16931 5952 16947 6016
rect 17011 5952 17017 6016
rect 16701 5951 17017 5952
rect 23003 6016 23319 6017
rect 23003 5952 23009 6016
rect 23073 5952 23089 6016
rect 23153 5952 23169 6016
rect 23233 5952 23249 6016
rect 23313 5952 23319 6016
rect 23003 5951 23319 5952
rect 20161 5674 20227 5677
rect 22553 5674 22619 5677
rect 20161 5672 22619 5674
rect 20161 5616 20166 5672
rect 20222 5616 22558 5672
rect 22614 5616 22619 5672
rect 20161 5614 22619 5616
rect 20161 5611 20227 5614
rect 22553 5611 22619 5614
rect 4757 5472 5073 5473
rect 4757 5408 4763 5472
rect 4827 5408 4843 5472
rect 4907 5408 4923 5472
rect 4987 5408 5003 5472
rect 5067 5408 5073 5472
rect 4757 5407 5073 5408
rect 11059 5472 11375 5473
rect 11059 5408 11065 5472
rect 11129 5408 11145 5472
rect 11209 5408 11225 5472
rect 11289 5408 11305 5472
rect 11369 5408 11375 5472
rect 11059 5407 11375 5408
rect 17361 5472 17677 5473
rect 17361 5408 17367 5472
rect 17431 5408 17447 5472
rect 17511 5408 17527 5472
rect 17591 5408 17607 5472
rect 17671 5408 17677 5472
rect 17361 5407 17677 5408
rect 23663 5472 23979 5473
rect 23663 5408 23669 5472
rect 23733 5408 23749 5472
rect 23813 5408 23829 5472
rect 23893 5408 23909 5472
rect 23973 5408 23979 5472
rect 23663 5407 23979 5408
rect 17125 5266 17191 5269
rect 17401 5266 17467 5269
rect 17125 5264 17467 5266
rect 17125 5208 17130 5264
rect 17186 5208 17406 5264
rect 17462 5208 17467 5264
rect 17125 5206 17467 5208
rect 17125 5203 17191 5206
rect 17401 5203 17467 5206
rect 4097 4928 4413 4929
rect 4097 4864 4103 4928
rect 4167 4864 4183 4928
rect 4247 4864 4263 4928
rect 4327 4864 4343 4928
rect 4407 4864 4413 4928
rect 4097 4863 4413 4864
rect 10399 4928 10715 4929
rect 10399 4864 10405 4928
rect 10469 4864 10485 4928
rect 10549 4864 10565 4928
rect 10629 4864 10645 4928
rect 10709 4864 10715 4928
rect 10399 4863 10715 4864
rect 16701 4928 17017 4929
rect 16701 4864 16707 4928
rect 16771 4864 16787 4928
rect 16851 4864 16867 4928
rect 16931 4864 16947 4928
rect 17011 4864 17017 4928
rect 16701 4863 17017 4864
rect 23003 4928 23319 4929
rect 23003 4864 23009 4928
rect 23073 4864 23089 4928
rect 23153 4864 23169 4928
rect 23233 4864 23249 4928
rect 23313 4864 23319 4928
rect 23003 4863 23319 4864
rect 13905 4586 13971 4589
rect 15285 4586 15351 4589
rect 13905 4584 15351 4586
rect 13905 4528 13910 4584
rect 13966 4528 15290 4584
rect 15346 4528 15351 4584
rect 13905 4526 15351 4528
rect 13905 4523 13971 4526
rect 15285 4523 15351 4526
rect 4757 4384 5073 4385
rect 4757 4320 4763 4384
rect 4827 4320 4843 4384
rect 4907 4320 4923 4384
rect 4987 4320 5003 4384
rect 5067 4320 5073 4384
rect 4757 4319 5073 4320
rect 11059 4384 11375 4385
rect 11059 4320 11065 4384
rect 11129 4320 11145 4384
rect 11209 4320 11225 4384
rect 11289 4320 11305 4384
rect 11369 4320 11375 4384
rect 11059 4319 11375 4320
rect 17361 4384 17677 4385
rect 17361 4320 17367 4384
rect 17431 4320 17447 4384
rect 17511 4320 17527 4384
rect 17591 4320 17607 4384
rect 17671 4320 17677 4384
rect 17361 4319 17677 4320
rect 23663 4384 23979 4385
rect 23663 4320 23669 4384
rect 23733 4320 23749 4384
rect 23813 4320 23829 4384
rect 23893 4320 23909 4384
rect 23973 4320 23979 4384
rect 23663 4319 23979 4320
rect 0 4178 800 4208
rect 3693 4178 3759 4181
rect 0 4176 3759 4178
rect 0 4120 3698 4176
rect 3754 4120 3759 4176
rect 0 4118 3759 4120
rect 0 4088 800 4118
rect 3693 4115 3759 4118
rect 25773 4178 25839 4181
rect 26681 4178 27481 4208
rect 25773 4176 27481 4178
rect 25773 4120 25778 4176
rect 25834 4120 27481 4176
rect 25773 4118 27481 4120
rect 25773 4115 25839 4118
rect 26681 4088 27481 4118
rect 4097 3840 4413 3841
rect 4097 3776 4103 3840
rect 4167 3776 4183 3840
rect 4247 3776 4263 3840
rect 4327 3776 4343 3840
rect 4407 3776 4413 3840
rect 4097 3775 4413 3776
rect 10399 3840 10715 3841
rect 10399 3776 10405 3840
rect 10469 3776 10485 3840
rect 10549 3776 10565 3840
rect 10629 3776 10645 3840
rect 10709 3776 10715 3840
rect 10399 3775 10715 3776
rect 16701 3840 17017 3841
rect 16701 3776 16707 3840
rect 16771 3776 16787 3840
rect 16851 3776 16867 3840
rect 16931 3776 16947 3840
rect 17011 3776 17017 3840
rect 16701 3775 17017 3776
rect 23003 3840 23319 3841
rect 23003 3776 23009 3840
rect 23073 3776 23089 3840
rect 23153 3776 23169 3840
rect 23233 3776 23249 3840
rect 23313 3776 23319 3840
rect 23003 3775 23319 3776
rect 4889 3498 4955 3501
rect 7465 3498 7531 3501
rect 4889 3496 7531 3498
rect 4889 3440 4894 3496
rect 4950 3440 7470 3496
rect 7526 3440 7531 3496
rect 4889 3438 7531 3440
rect 4889 3435 4955 3438
rect 7465 3435 7531 3438
rect 4757 3296 5073 3297
rect 4757 3232 4763 3296
rect 4827 3232 4843 3296
rect 4907 3232 4923 3296
rect 4987 3232 5003 3296
rect 5067 3232 5073 3296
rect 4757 3231 5073 3232
rect 11059 3296 11375 3297
rect 11059 3232 11065 3296
rect 11129 3232 11145 3296
rect 11209 3232 11225 3296
rect 11289 3232 11305 3296
rect 11369 3232 11375 3296
rect 11059 3231 11375 3232
rect 17361 3296 17677 3297
rect 17361 3232 17367 3296
rect 17431 3232 17447 3296
rect 17511 3232 17527 3296
rect 17591 3232 17607 3296
rect 17671 3232 17677 3296
rect 17361 3231 17677 3232
rect 23663 3296 23979 3297
rect 23663 3232 23669 3296
rect 23733 3232 23749 3296
rect 23813 3232 23829 3296
rect 23893 3232 23909 3296
rect 23973 3232 23979 3296
rect 23663 3231 23979 3232
rect 4097 2752 4413 2753
rect 4097 2688 4103 2752
rect 4167 2688 4183 2752
rect 4247 2688 4263 2752
rect 4327 2688 4343 2752
rect 4407 2688 4413 2752
rect 4097 2687 4413 2688
rect 10399 2752 10715 2753
rect 10399 2688 10405 2752
rect 10469 2688 10485 2752
rect 10549 2688 10565 2752
rect 10629 2688 10645 2752
rect 10709 2688 10715 2752
rect 10399 2687 10715 2688
rect 16701 2752 17017 2753
rect 16701 2688 16707 2752
rect 16771 2688 16787 2752
rect 16851 2688 16867 2752
rect 16931 2688 16947 2752
rect 17011 2688 17017 2752
rect 16701 2687 17017 2688
rect 23003 2752 23319 2753
rect 23003 2688 23009 2752
rect 23073 2688 23089 2752
rect 23153 2688 23169 2752
rect 23233 2688 23249 2752
rect 23313 2688 23319 2752
rect 23003 2687 23319 2688
rect 4757 2208 5073 2209
rect 4757 2144 4763 2208
rect 4827 2144 4843 2208
rect 4907 2144 4923 2208
rect 4987 2144 5003 2208
rect 5067 2144 5073 2208
rect 4757 2143 5073 2144
rect 11059 2208 11375 2209
rect 11059 2144 11065 2208
rect 11129 2144 11145 2208
rect 11209 2144 11225 2208
rect 11289 2144 11305 2208
rect 11369 2144 11375 2208
rect 11059 2143 11375 2144
rect 17361 2208 17677 2209
rect 17361 2144 17367 2208
rect 17431 2144 17447 2208
rect 17511 2144 17527 2208
rect 17591 2144 17607 2208
rect 17671 2144 17677 2208
rect 17361 2143 17677 2144
rect 23663 2208 23979 2209
rect 23663 2144 23669 2208
rect 23733 2144 23749 2208
rect 23813 2144 23829 2208
rect 23893 2144 23909 2208
rect 23973 2144 23979 2208
rect 23663 2143 23979 2144
rect 24761 98 24827 101
rect 26681 98 27481 128
rect 24761 96 27481 98
rect 24761 40 24766 96
rect 24822 40 27481 96
rect 24761 38 27481 40
rect 24761 35 24827 38
rect 26681 8 27481 38
<< via3 >>
rect 4763 27228 4827 27232
rect 4763 27172 4767 27228
rect 4767 27172 4823 27228
rect 4823 27172 4827 27228
rect 4763 27168 4827 27172
rect 4843 27228 4907 27232
rect 4843 27172 4847 27228
rect 4847 27172 4903 27228
rect 4903 27172 4907 27228
rect 4843 27168 4907 27172
rect 4923 27228 4987 27232
rect 4923 27172 4927 27228
rect 4927 27172 4983 27228
rect 4983 27172 4987 27228
rect 4923 27168 4987 27172
rect 5003 27228 5067 27232
rect 5003 27172 5007 27228
rect 5007 27172 5063 27228
rect 5063 27172 5067 27228
rect 5003 27168 5067 27172
rect 11065 27228 11129 27232
rect 11065 27172 11069 27228
rect 11069 27172 11125 27228
rect 11125 27172 11129 27228
rect 11065 27168 11129 27172
rect 11145 27228 11209 27232
rect 11145 27172 11149 27228
rect 11149 27172 11205 27228
rect 11205 27172 11209 27228
rect 11145 27168 11209 27172
rect 11225 27228 11289 27232
rect 11225 27172 11229 27228
rect 11229 27172 11285 27228
rect 11285 27172 11289 27228
rect 11225 27168 11289 27172
rect 11305 27228 11369 27232
rect 11305 27172 11309 27228
rect 11309 27172 11365 27228
rect 11365 27172 11369 27228
rect 11305 27168 11369 27172
rect 17367 27228 17431 27232
rect 17367 27172 17371 27228
rect 17371 27172 17427 27228
rect 17427 27172 17431 27228
rect 17367 27168 17431 27172
rect 17447 27228 17511 27232
rect 17447 27172 17451 27228
rect 17451 27172 17507 27228
rect 17507 27172 17511 27228
rect 17447 27168 17511 27172
rect 17527 27228 17591 27232
rect 17527 27172 17531 27228
rect 17531 27172 17587 27228
rect 17587 27172 17591 27228
rect 17527 27168 17591 27172
rect 17607 27228 17671 27232
rect 17607 27172 17611 27228
rect 17611 27172 17667 27228
rect 17667 27172 17671 27228
rect 17607 27168 17671 27172
rect 23669 27228 23733 27232
rect 23669 27172 23673 27228
rect 23673 27172 23729 27228
rect 23729 27172 23733 27228
rect 23669 27168 23733 27172
rect 23749 27228 23813 27232
rect 23749 27172 23753 27228
rect 23753 27172 23809 27228
rect 23809 27172 23813 27228
rect 23749 27168 23813 27172
rect 23829 27228 23893 27232
rect 23829 27172 23833 27228
rect 23833 27172 23889 27228
rect 23889 27172 23893 27228
rect 23829 27168 23893 27172
rect 23909 27228 23973 27232
rect 23909 27172 23913 27228
rect 23913 27172 23969 27228
rect 23969 27172 23973 27228
rect 23909 27168 23973 27172
rect 4103 26684 4167 26688
rect 4103 26628 4107 26684
rect 4107 26628 4163 26684
rect 4163 26628 4167 26684
rect 4103 26624 4167 26628
rect 4183 26684 4247 26688
rect 4183 26628 4187 26684
rect 4187 26628 4243 26684
rect 4243 26628 4247 26684
rect 4183 26624 4247 26628
rect 4263 26684 4327 26688
rect 4263 26628 4267 26684
rect 4267 26628 4323 26684
rect 4323 26628 4327 26684
rect 4263 26624 4327 26628
rect 4343 26684 4407 26688
rect 4343 26628 4347 26684
rect 4347 26628 4403 26684
rect 4403 26628 4407 26684
rect 4343 26624 4407 26628
rect 10405 26684 10469 26688
rect 10405 26628 10409 26684
rect 10409 26628 10465 26684
rect 10465 26628 10469 26684
rect 10405 26624 10469 26628
rect 10485 26684 10549 26688
rect 10485 26628 10489 26684
rect 10489 26628 10545 26684
rect 10545 26628 10549 26684
rect 10485 26624 10549 26628
rect 10565 26684 10629 26688
rect 10565 26628 10569 26684
rect 10569 26628 10625 26684
rect 10625 26628 10629 26684
rect 10565 26624 10629 26628
rect 10645 26684 10709 26688
rect 10645 26628 10649 26684
rect 10649 26628 10705 26684
rect 10705 26628 10709 26684
rect 10645 26624 10709 26628
rect 16707 26684 16771 26688
rect 16707 26628 16711 26684
rect 16711 26628 16767 26684
rect 16767 26628 16771 26684
rect 16707 26624 16771 26628
rect 16787 26684 16851 26688
rect 16787 26628 16791 26684
rect 16791 26628 16847 26684
rect 16847 26628 16851 26684
rect 16787 26624 16851 26628
rect 16867 26684 16931 26688
rect 16867 26628 16871 26684
rect 16871 26628 16927 26684
rect 16927 26628 16931 26684
rect 16867 26624 16931 26628
rect 16947 26684 17011 26688
rect 16947 26628 16951 26684
rect 16951 26628 17007 26684
rect 17007 26628 17011 26684
rect 16947 26624 17011 26628
rect 23009 26684 23073 26688
rect 23009 26628 23013 26684
rect 23013 26628 23069 26684
rect 23069 26628 23073 26684
rect 23009 26624 23073 26628
rect 23089 26684 23153 26688
rect 23089 26628 23093 26684
rect 23093 26628 23149 26684
rect 23149 26628 23153 26684
rect 23089 26624 23153 26628
rect 23169 26684 23233 26688
rect 23169 26628 23173 26684
rect 23173 26628 23229 26684
rect 23229 26628 23233 26684
rect 23169 26624 23233 26628
rect 23249 26684 23313 26688
rect 23249 26628 23253 26684
rect 23253 26628 23309 26684
rect 23309 26628 23313 26684
rect 23249 26624 23313 26628
rect 4763 26140 4827 26144
rect 4763 26084 4767 26140
rect 4767 26084 4823 26140
rect 4823 26084 4827 26140
rect 4763 26080 4827 26084
rect 4843 26140 4907 26144
rect 4843 26084 4847 26140
rect 4847 26084 4903 26140
rect 4903 26084 4907 26140
rect 4843 26080 4907 26084
rect 4923 26140 4987 26144
rect 4923 26084 4927 26140
rect 4927 26084 4983 26140
rect 4983 26084 4987 26140
rect 4923 26080 4987 26084
rect 5003 26140 5067 26144
rect 5003 26084 5007 26140
rect 5007 26084 5063 26140
rect 5063 26084 5067 26140
rect 5003 26080 5067 26084
rect 11065 26140 11129 26144
rect 11065 26084 11069 26140
rect 11069 26084 11125 26140
rect 11125 26084 11129 26140
rect 11065 26080 11129 26084
rect 11145 26140 11209 26144
rect 11145 26084 11149 26140
rect 11149 26084 11205 26140
rect 11205 26084 11209 26140
rect 11145 26080 11209 26084
rect 11225 26140 11289 26144
rect 11225 26084 11229 26140
rect 11229 26084 11285 26140
rect 11285 26084 11289 26140
rect 11225 26080 11289 26084
rect 11305 26140 11369 26144
rect 11305 26084 11309 26140
rect 11309 26084 11365 26140
rect 11365 26084 11369 26140
rect 11305 26080 11369 26084
rect 17367 26140 17431 26144
rect 17367 26084 17371 26140
rect 17371 26084 17427 26140
rect 17427 26084 17431 26140
rect 17367 26080 17431 26084
rect 17447 26140 17511 26144
rect 17447 26084 17451 26140
rect 17451 26084 17507 26140
rect 17507 26084 17511 26140
rect 17447 26080 17511 26084
rect 17527 26140 17591 26144
rect 17527 26084 17531 26140
rect 17531 26084 17587 26140
rect 17587 26084 17591 26140
rect 17527 26080 17591 26084
rect 17607 26140 17671 26144
rect 17607 26084 17611 26140
rect 17611 26084 17667 26140
rect 17667 26084 17671 26140
rect 17607 26080 17671 26084
rect 23669 26140 23733 26144
rect 23669 26084 23673 26140
rect 23673 26084 23729 26140
rect 23729 26084 23733 26140
rect 23669 26080 23733 26084
rect 23749 26140 23813 26144
rect 23749 26084 23753 26140
rect 23753 26084 23809 26140
rect 23809 26084 23813 26140
rect 23749 26080 23813 26084
rect 23829 26140 23893 26144
rect 23829 26084 23833 26140
rect 23833 26084 23889 26140
rect 23889 26084 23893 26140
rect 23829 26080 23893 26084
rect 23909 26140 23973 26144
rect 23909 26084 23913 26140
rect 23913 26084 23969 26140
rect 23969 26084 23973 26140
rect 23909 26080 23973 26084
rect 4103 25596 4167 25600
rect 4103 25540 4107 25596
rect 4107 25540 4163 25596
rect 4163 25540 4167 25596
rect 4103 25536 4167 25540
rect 4183 25596 4247 25600
rect 4183 25540 4187 25596
rect 4187 25540 4243 25596
rect 4243 25540 4247 25596
rect 4183 25536 4247 25540
rect 4263 25596 4327 25600
rect 4263 25540 4267 25596
rect 4267 25540 4323 25596
rect 4323 25540 4327 25596
rect 4263 25536 4327 25540
rect 4343 25596 4407 25600
rect 4343 25540 4347 25596
rect 4347 25540 4403 25596
rect 4403 25540 4407 25596
rect 4343 25536 4407 25540
rect 10405 25596 10469 25600
rect 10405 25540 10409 25596
rect 10409 25540 10465 25596
rect 10465 25540 10469 25596
rect 10405 25536 10469 25540
rect 10485 25596 10549 25600
rect 10485 25540 10489 25596
rect 10489 25540 10545 25596
rect 10545 25540 10549 25596
rect 10485 25536 10549 25540
rect 10565 25596 10629 25600
rect 10565 25540 10569 25596
rect 10569 25540 10625 25596
rect 10625 25540 10629 25596
rect 10565 25536 10629 25540
rect 10645 25596 10709 25600
rect 10645 25540 10649 25596
rect 10649 25540 10705 25596
rect 10705 25540 10709 25596
rect 10645 25536 10709 25540
rect 16707 25596 16771 25600
rect 16707 25540 16711 25596
rect 16711 25540 16767 25596
rect 16767 25540 16771 25596
rect 16707 25536 16771 25540
rect 16787 25596 16851 25600
rect 16787 25540 16791 25596
rect 16791 25540 16847 25596
rect 16847 25540 16851 25596
rect 16787 25536 16851 25540
rect 16867 25596 16931 25600
rect 16867 25540 16871 25596
rect 16871 25540 16927 25596
rect 16927 25540 16931 25596
rect 16867 25536 16931 25540
rect 16947 25596 17011 25600
rect 16947 25540 16951 25596
rect 16951 25540 17007 25596
rect 17007 25540 17011 25596
rect 16947 25536 17011 25540
rect 23009 25596 23073 25600
rect 23009 25540 23013 25596
rect 23013 25540 23069 25596
rect 23069 25540 23073 25596
rect 23009 25536 23073 25540
rect 23089 25596 23153 25600
rect 23089 25540 23093 25596
rect 23093 25540 23149 25596
rect 23149 25540 23153 25596
rect 23089 25536 23153 25540
rect 23169 25596 23233 25600
rect 23169 25540 23173 25596
rect 23173 25540 23229 25596
rect 23229 25540 23233 25596
rect 23169 25536 23233 25540
rect 23249 25596 23313 25600
rect 23249 25540 23253 25596
rect 23253 25540 23309 25596
rect 23309 25540 23313 25596
rect 23249 25536 23313 25540
rect 4763 25052 4827 25056
rect 4763 24996 4767 25052
rect 4767 24996 4823 25052
rect 4823 24996 4827 25052
rect 4763 24992 4827 24996
rect 4843 25052 4907 25056
rect 4843 24996 4847 25052
rect 4847 24996 4903 25052
rect 4903 24996 4907 25052
rect 4843 24992 4907 24996
rect 4923 25052 4987 25056
rect 4923 24996 4927 25052
rect 4927 24996 4983 25052
rect 4983 24996 4987 25052
rect 4923 24992 4987 24996
rect 5003 25052 5067 25056
rect 5003 24996 5007 25052
rect 5007 24996 5063 25052
rect 5063 24996 5067 25052
rect 5003 24992 5067 24996
rect 11065 25052 11129 25056
rect 11065 24996 11069 25052
rect 11069 24996 11125 25052
rect 11125 24996 11129 25052
rect 11065 24992 11129 24996
rect 11145 25052 11209 25056
rect 11145 24996 11149 25052
rect 11149 24996 11205 25052
rect 11205 24996 11209 25052
rect 11145 24992 11209 24996
rect 11225 25052 11289 25056
rect 11225 24996 11229 25052
rect 11229 24996 11285 25052
rect 11285 24996 11289 25052
rect 11225 24992 11289 24996
rect 11305 25052 11369 25056
rect 11305 24996 11309 25052
rect 11309 24996 11365 25052
rect 11365 24996 11369 25052
rect 11305 24992 11369 24996
rect 17367 25052 17431 25056
rect 17367 24996 17371 25052
rect 17371 24996 17427 25052
rect 17427 24996 17431 25052
rect 17367 24992 17431 24996
rect 17447 25052 17511 25056
rect 17447 24996 17451 25052
rect 17451 24996 17507 25052
rect 17507 24996 17511 25052
rect 17447 24992 17511 24996
rect 17527 25052 17591 25056
rect 17527 24996 17531 25052
rect 17531 24996 17587 25052
rect 17587 24996 17591 25052
rect 17527 24992 17591 24996
rect 17607 25052 17671 25056
rect 17607 24996 17611 25052
rect 17611 24996 17667 25052
rect 17667 24996 17671 25052
rect 17607 24992 17671 24996
rect 23669 25052 23733 25056
rect 23669 24996 23673 25052
rect 23673 24996 23729 25052
rect 23729 24996 23733 25052
rect 23669 24992 23733 24996
rect 23749 25052 23813 25056
rect 23749 24996 23753 25052
rect 23753 24996 23809 25052
rect 23809 24996 23813 25052
rect 23749 24992 23813 24996
rect 23829 25052 23893 25056
rect 23829 24996 23833 25052
rect 23833 24996 23889 25052
rect 23889 24996 23893 25052
rect 23829 24992 23893 24996
rect 23909 25052 23973 25056
rect 23909 24996 23913 25052
rect 23913 24996 23969 25052
rect 23969 24996 23973 25052
rect 23909 24992 23973 24996
rect 4103 24508 4167 24512
rect 4103 24452 4107 24508
rect 4107 24452 4163 24508
rect 4163 24452 4167 24508
rect 4103 24448 4167 24452
rect 4183 24508 4247 24512
rect 4183 24452 4187 24508
rect 4187 24452 4243 24508
rect 4243 24452 4247 24508
rect 4183 24448 4247 24452
rect 4263 24508 4327 24512
rect 4263 24452 4267 24508
rect 4267 24452 4323 24508
rect 4323 24452 4327 24508
rect 4263 24448 4327 24452
rect 4343 24508 4407 24512
rect 4343 24452 4347 24508
rect 4347 24452 4403 24508
rect 4403 24452 4407 24508
rect 4343 24448 4407 24452
rect 10405 24508 10469 24512
rect 10405 24452 10409 24508
rect 10409 24452 10465 24508
rect 10465 24452 10469 24508
rect 10405 24448 10469 24452
rect 10485 24508 10549 24512
rect 10485 24452 10489 24508
rect 10489 24452 10545 24508
rect 10545 24452 10549 24508
rect 10485 24448 10549 24452
rect 10565 24508 10629 24512
rect 10565 24452 10569 24508
rect 10569 24452 10625 24508
rect 10625 24452 10629 24508
rect 10565 24448 10629 24452
rect 10645 24508 10709 24512
rect 10645 24452 10649 24508
rect 10649 24452 10705 24508
rect 10705 24452 10709 24508
rect 10645 24448 10709 24452
rect 16707 24508 16771 24512
rect 16707 24452 16711 24508
rect 16711 24452 16767 24508
rect 16767 24452 16771 24508
rect 16707 24448 16771 24452
rect 16787 24508 16851 24512
rect 16787 24452 16791 24508
rect 16791 24452 16847 24508
rect 16847 24452 16851 24508
rect 16787 24448 16851 24452
rect 16867 24508 16931 24512
rect 16867 24452 16871 24508
rect 16871 24452 16927 24508
rect 16927 24452 16931 24508
rect 16867 24448 16931 24452
rect 16947 24508 17011 24512
rect 16947 24452 16951 24508
rect 16951 24452 17007 24508
rect 17007 24452 17011 24508
rect 16947 24448 17011 24452
rect 23009 24508 23073 24512
rect 23009 24452 23013 24508
rect 23013 24452 23069 24508
rect 23069 24452 23073 24508
rect 23009 24448 23073 24452
rect 23089 24508 23153 24512
rect 23089 24452 23093 24508
rect 23093 24452 23149 24508
rect 23149 24452 23153 24508
rect 23089 24448 23153 24452
rect 23169 24508 23233 24512
rect 23169 24452 23173 24508
rect 23173 24452 23229 24508
rect 23229 24452 23233 24508
rect 23169 24448 23233 24452
rect 23249 24508 23313 24512
rect 23249 24452 23253 24508
rect 23253 24452 23309 24508
rect 23309 24452 23313 24508
rect 23249 24448 23313 24452
rect 4763 23964 4827 23968
rect 4763 23908 4767 23964
rect 4767 23908 4823 23964
rect 4823 23908 4827 23964
rect 4763 23904 4827 23908
rect 4843 23964 4907 23968
rect 4843 23908 4847 23964
rect 4847 23908 4903 23964
rect 4903 23908 4907 23964
rect 4843 23904 4907 23908
rect 4923 23964 4987 23968
rect 4923 23908 4927 23964
rect 4927 23908 4983 23964
rect 4983 23908 4987 23964
rect 4923 23904 4987 23908
rect 5003 23964 5067 23968
rect 5003 23908 5007 23964
rect 5007 23908 5063 23964
rect 5063 23908 5067 23964
rect 5003 23904 5067 23908
rect 11065 23964 11129 23968
rect 11065 23908 11069 23964
rect 11069 23908 11125 23964
rect 11125 23908 11129 23964
rect 11065 23904 11129 23908
rect 11145 23964 11209 23968
rect 11145 23908 11149 23964
rect 11149 23908 11205 23964
rect 11205 23908 11209 23964
rect 11145 23904 11209 23908
rect 11225 23964 11289 23968
rect 11225 23908 11229 23964
rect 11229 23908 11285 23964
rect 11285 23908 11289 23964
rect 11225 23904 11289 23908
rect 11305 23964 11369 23968
rect 11305 23908 11309 23964
rect 11309 23908 11365 23964
rect 11365 23908 11369 23964
rect 11305 23904 11369 23908
rect 17367 23964 17431 23968
rect 17367 23908 17371 23964
rect 17371 23908 17427 23964
rect 17427 23908 17431 23964
rect 17367 23904 17431 23908
rect 17447 23964 17511 23968
rect 17447 23908 17451 23964
rect 17451 23908 17507 23964
rect 17507 23908 17511 23964
rect 17447 23904 17511 23908
rect 17527 23964 17591 23968
rect 17527 23908 17531 23964
rect 17531 23908 17587 23964
rect 17587 23908 17591 23964
rect 17527 23904 17591 23908
rect 17607 23964 17671 23968
rect 17607 23908 17611 23964
rect 17611 23908 17667 23964
rect 17667 23908 17671 23964
rect 17607 23904 17671 23908
rect 23669 23964 23733 23968
rect 23669 23908 23673 23964
rect 23673 23908 23729 23964
rect 23729 23908 23733 23964
rect 23669 23904 23733 23908
rect 23749 23964 23813 23968
rect 23749 23908 23753 23964
rect 23753 23908 23809 23964
rect 23809 23908 23813 23964
rect 23749 23904 23813 23908
rect 23829 23964 23893 23968
rect 23829 23908 23833 23964
rect 23833 23908 23889 23964
rect 23889 23908 23893 23964
rect 23829 23904 23893 23908
rect 23909 23964 23973 23968
rect 23909 23908 23913 23964
rect 23913 23908 23969 23964
rect 23969 23908 23973 23964
rect 23909 23904 23973 23908
rect 5580 23488 5644 23492
rect 5580 23432 5594 23488
rect 5594 23432 5644 23488
rect 5580 23428 5644 23432
rect 4103 23420 4167 23424
rect 4103 23364 4107 23420
rect 4107 23364 4163 23420
rect 4163 23364 4167 23420
rect 4103 23360 4167 23364
rect 4183 23420 4247 23424
rect 4183 23364 4187 23420
rect 4187 23364 4243 23420
rect 4243 23364 4247 23420
rect 4183 23360 4247 23364
rect 4263 23420 4327 23424
rect 4263 23364 4267 23420
rect 4267 23364 4323 23420
rect 4323 23364 4327 23420
rect 4263 23360 4327 23364
rect 4343 23420 4407 23424
rect 4343 23364 4347 23420
rect 4347 23364 4403 23420
rect 4403 23364 4407 23420
rect 4343 23360 4407 23364
rect 10405 23420 10469 23424
rect 10405 23364 10409 23420
rect 10409 23364 10465 23420
rect 10465 23364 10469 23420
rect 10405 23360 10469 23364
rect 10485 23420 10549 23424
rect 10485 23364 10489 23420
rect 10489 23364 10545 23420
rect 10545 23364 10549 23420
rect 10485 23360 10549 23364
rect 10565 23420 10629 23424
rect 10565 23364 10569 23420
rect 10569 23364 10625 23420
rect 10625 23364 10629 23420
rect 10565 23360 10629 23364
rect 10645 23420 10709 23424
rect 10645 23364 10649 23420
rect 10649 23364 10705 23420
rect 10705 23364 10709 23420
rect 10645 23360 10709 23364
rect 16707 23420 16771 23424
rect 16707 23364 16711 23420
rect 16711 23364 16767 23420
rect 16767 23364 16771 23420
rect 16707 23360 16771 23364
rect 16787 23420 16851 23424
rect 16787 23364 16791 23420
rect 16791 23364 16847 23420
rect 16847 23364 16851 23420
rect 16787 23360 16851 23364
rect 16867 23420 16931 23424
rect 16867 23364 16871 23420
rect 16871 23364 16927 23420
rect 16927 23364 16931 23420
rect 16867 23360 16931 23364
rect 16947 23420 17011 23424
rect 16947 23364 16951 23420
rect 16951 23364 17007 23420
rect 17007 23364 17011 23420
rect 16947 23360 17011 23364
rect 23009 23420 23073 23424
rect 23009 23364 23013 23420
rect 23013 23364 23069 23420
rect 23069 23364 23073 23420
rect 23009 23360 23073 23364
rect 23089 23420 23153 23424
rect 23089 23364 23093 23420
rect 23093 23364 23149 23420
rect 23149 23364 23153 23420
rect 23089 23360 23153 23364
rect 23169 23420 23233 23424
rect 23169 23364 23173 23420
rect 23173 23364 23229 23420
rect 23229 23364 23233 23420
rect 23169 23360 23233 23364
rect 23249 23420 23313 23424
rect 23249 23364 23253 23420
rect 23253 23364 23309 23420
rect 23309 23364 23313 23420
rect 23249 23360 23313 23364
rect 4763 22876 4827 22880
rect 4763 22820 4767 22876
rect 4767 22820 4823 22876
rect 4823 22820 4827 22876
rect 4763 22816 4827 22820
rect 4843 22876 4907 22880
rect 4843 22820 4847 22876
rect 4847 22820 4903 22876
rect 4903 22820 4907 22876
rect 4843 22816 4907 22820
rect 4923 22876 4987 22880
rect 4923 22820 4927 22876
rect 4927 22820 4983 22876
rect 4983 22820 4987 22876
rect 4923 22816 4987 22820
rect 5003 22876 5067 22880
rect 5003 22820 5007 22876
rect 5007 22820 5063 22876
rect 5063 22820 5067 22876
rect 5003 22816 5067 22820
rect 11065 22876 11129 22880
rect 11065 22820 11069 22876
rect 11069 22820 11125 22876
rect 11125 22820 11129 22876
rect 11065 22816 11129 22820
rect 11145 22876 11209 22880
rect 11145 22820 11149 22876
rect 11149 22820 11205 22876
rect 11205 22820 11209 22876
rect 11145 22816 11209 22820
rect 11225 22876 11289 22880
rect 11225 22820 11229 22876
rect 11229 22820 11285 22876
rect 11285 22820 11289 22876
rect 11225 22816 11289 22820
rect 11305 22876 11369 22880
rect 11305 22820 11309 22876
rect 11309 22820 11365 22876
rect 11365 22820 11369 22876
rect 11305 22816 11369 22820
rect 17367 22876 17431 22880
rect 17367 22820 17371 22876
rect 17371 22820 17427 22876
rect 17427 22820 17431 22876
rect 17367 22816 17431 22820
rect 17447 22876 17511 22880
rect 17447 22820 17451 22876
rect 17451 22820 17507 22876
rect 17507 22820 17511 22876
rect 17447 22816 17511 22820
rect 17527 22876 17591 22880
rect 17527 22820 17531 22876
rect 17531 22820 17587 22876
rect 17587 22820 17591 22876
rect 17527 22816 17591 22820
rect 17607 22876 17671 22880
rect 17607 22820 17611 22876
rect 17611 22820 17667 22876
rect 17667 22820 17671 22876
rect 17607 22816 17671 22820
rect 23669 22876 23733 22880
rect 23669 22820 23673 22876
rect 23673 22820 23729 22876
rect 23729 22820 23733 22876
rect 23669 22816 23733 22820
rect 23749 22876 23813 22880
rect 23749 22820 23753 22876
rect 23753 22820 23809 22876
rect 23809 22820 23813 22876
rect 23749 22816 23813 22820
rect 23829 22876 23893 22880
rect 23829 22820 23833 22876
rect 23833 22820 23889 22876
rect 23889 22820 23893 22876
rect 23829 22816 23893 22820
rect 23909 22876 23973 22880
rect 23909 22820 23913 22876
rect 23913 22820 23969 22876
rect 23969 22820 23973 22876
rect 23909 22816 23973 22820
rect 4103 22332 4167 22336
rect 4103 22276 4107 22332
rect 4107 22276 4163 22332
rect 4163 22276 4167 22332
rect 4103 22272 4167 22276
rect 4183 22332 4247 22336
rect 4183 22276 4187 22332
rect 4187 22276 4243 22332
rect 4243 22276 4247 22332
rect 4183 22272 4247 22276
rect 4263 22332 4327 22336
rect 4263 22276 4267 22332
rect 4267 22276 4323 22332
rect 4323 22276 4327 22332
rect 4263 22272 4327 22276
rect 4343 22332 4407 22336
rect 4343 22276 4347 22332
rect 4347 22276 4403 22332
rect 4403 22276 4407 22332
rect 4343 22272 4407 22276
rect 10405 22332 10469 22336
rect 10405 22276 10409 22332
rect 10409 22276 10465 22332
rect 10465 22276 10469 22332
rect 10405 22272 10469 22276
rect 10485 22332 10549 22336
rect 10485 22276 10489 22332
rect 10489 22276 10545 22332
rect 10545 22276 10549 22332
rect 10485 22272 10549 22276
rect 10565 22332 10629 22336
rect 10565 22276 10569 22332
rect 10569 22276 10625 22332
rect 10625 22276 10629 22332
rect 10565 22272 10629 22276
rect 10645 22332 10709 22336
rect 10645 22276 10649 22332
rect 10649 22276 10705 22332
rect 10705 22276 10709 22332
rect 10645 22272 10709 22276
rect 16707 22332 16771 22336
rect 16707 22276 16711 22332
rect 16711 22276 16767 22332
rect 16767 22276 16771 22332
rect 16707 22272 16771 22276
rect 16787 22332 16851 22336
rect 16787 22276 16791 22332
rect 16791 22276 16847 22332
rect 16847 22276 16851 22332
rect 16787 22272 16851 22276
rect 16867 22332 16931 22336
rect 16867 22276 16871 22332
rect 16871 22276 16927 22332
rect 16927 22276 16931 22332
rect 16867 22272 16931 22276
rect 16947 22332 17011 22336
rect 16947 22276 16951 22332
rect 16951 22276 17007 22332
rect 17007 22276 17011 22332
rect 16947 22272 17011 22276
rect 23009 22332 23073 22336
rect 23009 22276 23013 22332
rect 23013 22276 23069 22332
rect 23069 22276 23073 22332
rect 23009 22272 23073 22276
rect 23089 22332 23153 22336
rect 23089 22276 23093 22332
rect 23093 22276 23149 22332
rect 23149 22276 23153 22332
rect 23089 22272 23153 22276
rect 23169 22332 23233 22336
rect 23169 22276 23173 22332
rect 23173 22276 23229 22332
rect 23229 22276 23233 22332
rect 23169 22272 23233 22276
rect 23249 22332 23313 22336
rect 23249 22276 23253 22332
rect 23253 22276 23309 22332
rect 23309 22276 23313 22332
rect 23249 22272 23313 22276
rect 6132 21932 6196 21996
rect 4763 21788 4827 21792
rect 4763 21732 4767 21788
rect 4767 21732 4823 21788
rect 4823 21732 4827 21788
rect 4763 21728 4827 21732
rect 4843 21788 4907 21792
rect 4843 21732 4847 21788
rect 4847 21732 4903 21788
rect 4903 21732 4907 21788
rect 4843 21728 4907 21732
rect 4923 21788 4987 21792
rect 4923 21732 4927 21788
rect 4927 21732 4983 21788
rect 4983 21732 4987 21788
rect 4923 21728 4987 21732
rect 5003 21788 5067 21792
rect 5003 21732 5007 21788
rect 5007 21732 5063 21788
rect 5063 21732 5067 21788
rect 5003 21728 5067 21732
rect 11065 21788 11129 21792
rect 11065 21732 11069 21788
rect 11069 21732 11125 21788
rect 11125 21732 11129 21788
rect 11065 21728 11129 21732
rect 11145 21788 11209 21792
rect 11145 21732 11149 21788
rect 11149 21732 11205 21788
rect 11205 21732 11209 21788
rect 11145 21728 11209 21732
rect 11225 21788 11289 21792
rect 11225 21732 11229 21788
rect 11229 21732 11285 21788
rect 11285 21732 11289 21788
rect 11225 21728 11289 21732
rect 11305 21788 11369 21792
rect 11305 21732 11309 21788
rect 11309 21732 11365 21788
rect 11365 21732 11369 21788
rect 11305 21728 11369 21732
rect 17367 21788 17431 21792
rect 17367 21732 17371 21788
rect 17371 21732 17427 21788
rect 17427 21732 17431 21788
rect 17367 21728 17431 21732
rect 17447 21788 17511 21792
rect 17447 21732 17451 21788
rect 17451 21732 17507 21788
rect 17507 21732 17511 21788
rect 17447 21728 17511 21732
rect 17527 21788 17591 21792
rect 17527 21732 17531 21788
rect 17531 21732 17587 21788
rect 17587 21732 17591 21788
rect 17527 21728 17591 21732
rect 17607 21788 17671 21792
rect 17607 21732 17611 21788
rect 17611 21732 17667 21788
rect 17667 21732 17671 21788
rect 17607 21728 17671 21732
rect 23669 21788 23733 21792
rect 23669 21732 23673 21788
rect 23673 21732 23729 21788
rect 23729 21732 23733 21788
rect 23669 21728 23733 21732
rect 23749 21788 23813 21792
rect 23749 21732 23753 21788
rect 23753 21732 23809 21788
rect 23809 21732 23813 21788
rect 23749 21728 23813 21732
rect 23829 21788 23893 21792
rect 23829 21732 23833 21788
rect 23833 21732 23889 21788
rect 23889 21732 23893 21788
rect 23829 21728 23893 21732
rect 23909 21788 23973 21792
rect 23909 21732 23913 21788
rect 23913 21732 23969 21788
rect 23969 21732 23973 21788
rect 23909 21728 23973 21732
rect 4103 21244 4167 21248
rect 4103 21188 4107 21244
rect 4107 21188 4163 21244
rect 4163 21188 4167 21244
rect 4103 21184 4167 21188
rect 4183 21244 4247 21248
rect 4183 21188 4187 21244
rect 4187 21188 4243 21244
rect 4243 21188 4247 21244
rect 4183 21184 4247 21188
rect 4263 21244 4327 21248
rect 4263 21188 4267 21244
rect 4267 21188 4323 21244
rect 4323 21188 4327 21244
rect 4263 21184 4327 21188
rect 4343 21244 4407 21248
rect 4343 21188 4347 21244
rect 4347 21188 4403 21244
rect 4403 21188 4407 21244
rect 4343 21184 4407 21188
rect 10405 21244 10469 21248
rect 10405 21188 10409 21244
rect 10409 21188 10465 21244
rect 10465 21188 10469 21244
rect 10405 21184 10469 21188
rect 10485 21244 10549 21248
rect 10485 21188 10489 21244
rect 10489 21188 10545 21244
rect 10545 21188 10549 21244
rect 10485 21184 10549 21188
rect 10565 21244 10629 21248
rect 10565 21188 10569 21244
rect 10569 21188 10625 21244
rect 10625 21188 10629 21244
rect 10565 21184 10629 21188
rect 10645 21244 10709 21248
rect 10645 21188 10649 21244
rect 10649 21188 10705 21244
rect 10705 21188 10709 21244
rect 10645 21184 10709 21188
rect 16707 21244 16771 21248
rect 16707 21188 16711 21244
rect 16711 21188 16767 21244
rect 16767 21188 16771 21244
rect 16707 21184 16771 21188
rect 16787 21244 16851 21248
rect 16787 21188 16791 21244
rect 16791 21188 16847 21244
rect 16847 21188 16851 21244
rect 16787 21184 16851 21188
rect 16867 21244 16931 21248
rect 16867 21188 16871 21244
rect 16871 21188 16927 21244
rect 16927 21188 16931 21244
rect 16867 21184 16931 21188
rect 16947 21244 17011 21248
rect 16947 21188 16951 21244
rect 16951 21188 17007 21244
rect 17007 21188 17011 21244
rect 16947 21184 17011 21188
rect 23009 21244 23073 21248
rect 23009 21188 23013 21244
rect 23013 21188 23069 21244
rect 23069 21188 23073 21244
rect 23009 21184 23073 21188
rect 23089 21244 23153 21248
rect 23089 21188 23093 21244
rect 23093 21188 23149 21244
rect 23149 21188 23153 21244
rect 23089 21184 23153 21188
rect 23169 21244 23233 21248
rect 23169 21188 23173 21244
rect 23173 21188 23229 21244
rect 23229 21188 23233 21244
rect 23169 21184 23233 21188
rect 23249 21244 23313 21248
rect 23249 21188 23253 21244
rect 23253 21188 23309 21244
rect 23309 21188 23313 21244
rect 23249 21184 23313 21188
rect 4763 20700 4827 20704
rect 4763 20644 4767 20700
rect 4767 20644 4823 20700
rect 4823 20644 4827 20700
rect 4763 20640 4827 20644
rect 4843 20700 4907 20704
rect 4843 20644 4847 20700
rect 4847 20644 4903 20700
rect 4903 20644 4907 20700
rect 4843 20640 4907 20644
rect 4923 20700 4987 20704
rect 4923 20644 4927 20700
rect 4927 20644 4983 20700
rect 4983 20644 4987 20700
rect 4923 20640 4987 20644
rect 5003 20700 5067 20704
rect 5003 20644 5007 20700
rect 5007 20644 5063 20700
rect 5063 20644 5067 20700
rect 5003 20640 5067 20644
rect 11065 20700 11129 20704
rect 11065 20644 11069 20700
rect 11069 20644 11125 20700
rect 11125 20644 11129 20700
rect 11065 20640 11129 20644
rect 11145 20700 11209 20704
rect 11145 20644 11149 20700
rect 11149 20644 11205 20700
rect 11205 20644 11209 20700
rect 11145 20640 11209 20644
rect 11225 20700 11289 20704
rect 11225 20644 11229 20700
rect 11229 20644 11285 20700
rect 11285 20644 11289 20700
rect 11225 20640 11289 20644
rect 11305 20700 11369 20704
rect 11305 20644 11309 20700
rect 11309 20644 11365 20700
rect 11365 20644 11369 20700
rect 11305 20640 11369 20644
rect 17367 20700 17431 20704
rect 17367 20644 17371 20700
rect 17371 20644 17427 20700
rect 17427 20644 17431 20700
rect 17367 20640 17431 20644
rect 17447 20700 17511 20704
rect 17447 20644 17451 20700
rect 17451 20644 17507 20700
rect 17507 20644 17511 20700
rect 17447 20640 17511 20644
rect 17527 20700 17591 20704
rect 17527 20644 17531 20700
rect 17531 20644 17587 20700
rect 17587 20644 17591 20700
rect 17527 20640 17591 20644
rect 17607 20700 17671 20704
rect 17607 20644 17611 20700
rect 17611 20644 17667 20700
rect 17667 20644 17671 20700
rect 17607 20640 17671 20644
rect 23669 20700 23733 20704
rect 23669 20644 23673 20700
rect 23673 20644 23729 20700
rect 23729 20644 23733 20700
rect 23669 20640 23733 20644
rect 23749 20700 23813 20704
rect 23749 20644 23753 20700
rect 23753 20644 23809 20700
rect 23809 20644 23813 20700
rect 23749 20640 23813 20644
rect 23829 20700 23893 20704
rect 23829 20644 23833 20700
rect 23833 20644 23889 20700
rect 23889 20644 23893 20700
rect 23829 20640 23893 20644
rect 23909 20700 23973 20704
rect 23909 20644 23913 20700
rect 23913 20644 23969 20700
rect 23969 20644 23973 20700
rect 23909 20640 23973 20644
rect 4103 20156 4167 20160
rect 4103 20100 4107 20156
rect 4107 20100 4163 20156
rect 4163 20100 4167 20156
rect 4103 20096 4167 20100
rect 4183 20156 4247 20160
rect 4183 20100 4187 20156
rect 4187 20100 4243 20156
rect 4243 20100 4247 20156
rect 4183 20096 4247 20100
rect 4263 20156 4327 20160
rect 4263 20100 4267 20156
rect 4267 20100 4323 20156
rect 4323 20100 4327 20156
rect 4263 20096 4327 20100
rect 4343 20156 4407 20160
rect 4343 20100 4347 20156
rect 4347 20100 4403 20156
rect 4403 20100 4407 20156
rect 4343 20096 4407 20100
rect 10405 20156 10469 20160
rect 10405 20100 10409 20156
rect 10409 20100 10465 20156
rect 10465 20100 10469 20156
rect 10405 20096 10469 20100
rect 10485 20156 10549 20160
rect 10485 20100 10489 20156
rect 10489 20100 10545 20156
rect 10545 20100 10549 20156
rect 10485 20096 10549 20100
rect 10565 20156 10629 20160
rect 10565 20100 10569 20156
rect 10569 20100 10625 20156
rect 10625 20100 10629 20156
rect 10565 20096 10629 20100
rect 10645 20156 10709 20160
rect 10645 20100 10649 20156
rect 10649 20100 10705 20156
rect 10705 20100 10709 20156
rect 10645 20096 10709 20100
rect 16707 20156 16771 20160
rect 16707 20100 16711 20156
rect 16711 20100 16767 20156
rect 16767 20100 16771 20156
rect 16707 20096 16771 20100
rect 16787 20156 16851 20160
rect 16787 20100 16791 20156
rect 16791 20100 16847 20156
rect 16847 20100 16851 20156
rect 16787 20096 16851 20100
rect 16867 20156 16931 20160
rect 16867 20100 16871 20156
rect 16871 20100 16927 20156
rect 16927 20100 16931 20156
rect 16867 20096 16931 20100
rect 16947 20156 17011 20160
rect 16947 20100 16951 20156
rect 16951 20100 17007 20156
rect 17007 20100 17011 20156
rect 16947 20096 17011 20100
rect 23009 20156 23073 20160
rect 23009 20100 23013 20156
rect 23013 20100 23069 20156
rect 23069 20100 23073 20156
rect 23009 20096 23073 20100
rect 23089 20156 23153 20160
rect 23089 20100 23093 20156
rect 23093 20100 23149 20156
rect 23149 20100 23153 20156
rect 23089 20096 23153 20100
rect 23169 20156 23233 20160
rect 23169 20100 23173 20156
rect 23173 20100 23229 20156
rect 23229 20100 23233 20156
rect 23169 20096 23233 20100
rect 23249 20156 23313 20160
rect 23249 20100 23253 20156
rect 23253 20100 23309 20156
rect 23309 20100 23313 20156
rect 23249 20096 23313 20100
rect 4763 19612 4827 19616
rect 4763 19556 4767 19612
rect 4767 19556 4823 19612
rect 4823 19556 4827 19612
rect 4763 19552 4827 19556
rect 4843 19612 4907 19616
rect 4843 19556 4847 19612
rect 4847 19556 4903 19612
rect 4903 19556 4907 19612
rect 4843 19552 4907 19556
rect 4923 19612 4987 19616
rect 4923 19556 4927 19612
rect 4927 19556 4983 19612
rect 4983 19556 4987 19612
rect 4923 19552 4987 19556
rect 5003 19612 5067 19616
rect 5003 19556 5007 19612
rect 5007 19556 5063 19612
rect 5063 19556 5067 19612
rect 5003 19552 5067 19556
rect 11065 19612 11129 19616
rect 11065 19556 11069 19612
rect 11069 19556 11125 19612
rect 11125 19556 11129 19612
rect 11065 19552 11129 19556
rect 11145 19612 11209 19616
rect 11145 19556 11149 19612
rect 11149 19556 11205 19612
rect 11205 19556 11209 19612
rect 11145 19552 11209 19556
rect 11225 19612 11289 19616
rect 11225 19556 11229 19612
rect 11229 19556 11285 19612
rect 11285 19556 11289 19612
rect 11225 19552 11289 19556
rect 11305 19612 11369 19616
rect 11305 19556 11309 19612
rect 11309 19556 11365 19612
rect 11365 19556 11369 19612
rect 11305 19552 11369 19556
rect 17367 19612 17431 19616
rect 17367 19556 17371 19612
rect 17371 19556 17427 19612
rect 17427 19556 17431 19612
rect 17367 19552 17431 19556
rect 17447 19612 17511 19616
rect 17447 19556 17451 19612
rect 17451 19556 17507 19612
rect 17507 19556 17511 19612
rect 17447 19552 17511 19556
rect 17527 19612 17591 19616
rect 17527 19556 17531 19612
rect 17531 19556 17587 19612
rect 17587 19556 17591 19612
rect 17527 19552 17591 19556
rect 17607 19612 17671 19616
rect 17607 19556 17611 19612
rect 17611 19556 17667 19612
rect 17667 19556 17671 19612
rect 17607 19552 17671 19556
rect 23669 19612 23733 19616
rect 23669 19556 23673 19612
rect 23673 19556 23729 19612
rect 23729 19556 23733 19612
rect 23669 19552 23733 19556
rect 23749 19612 23813 19616
rect 23749 19556 23753 19612
rect 23753 19556 23809 19612
rect 23809 19556 23813 19612
rect 23749 19552 23813 19556
rect 23829 19612 23893 19616
rect 23829 19556 23833 19612
rect 23833 19556 23889 19612
rect 23889 19556 23893 19612
rect 23829 19552 23893 19556
rect 23909 19612 23973 19616
rect 23909 19556 23913 19612
rect 23913 19556 23969 19612
rect 23969 19556 23973 19612
rect 23909 19552 23973 19556
rect 4103 19068 4167 19072
rect 4103 19012 4107 19068
rect 4107 19012 4163 19068
rect 4163 19012 4167 19068
rect 4103 19008 4167 19012
rect 4183 19068 4247 19072
rect 4183 19012 4187 19068
rect 4187 19012 4243 19068
rect 4243 19012 4247 19068
rect 4183 19008 4247 19012
rect 4263 19068 4327 19072
rect 4263 19012 4267 19068
rect 4267 19012 4323 19068
rect 4323 19012 4327 19068
rect 4263 19008 4327 19012
rect 4343 19068 4407 19072
rect 4343 19012 4347 19068
rect 4347 19012 4403 19068
rect 4403 19012 4407 19068
rect 4343 19008 4407 19012
rect 10405 19068 10469 19072
rect 10405 19012 10409 19068
rect 10409 19012 10465 19068
rect 10465 19012 10469 19068
rect 10405 19008 10469 19012
rect 10485 19068 10549 19072
rect 10485 19012 10489 19068
rect 10489 19012 10545 19068
rect 10545 19012 10549 19068
rect 10485 19008 10549 19012
rect 10565 19068 10629 19072
rect 10565 19012 10569 19068
rect 10569 19012 10625 19068
rect 10625 19012 10629 19068
rect 10565 19008 10629 19012
rect 10645 19068 10709 19072
rect 10645 19012 10649 19068
rect 10649 19012 10705 19068
rect 10705 19012 10709 19068
rect 10645 19008 10709 19012
rect 16707 19068 16771 19072
rect 16707 19012 16711 19068
rect 16711 19012 16767 19068
rect 16767 19012 16771 19068
rect 16707 19008 16771 19012
rect 16787 19068 16851 19072
rect 16787 19012 16791 19068
rect 16791 19012 16847 19068
rect 16847 19012 16851 19068
rect 16787 19008 16851 19012
rect 16867 19068 16931 19072
rect 16867 19012 16871 19068
rect 16871 19012 16927 19068
rect 16927 19012 16931 19068
rect 16867 19008 16931 19012
rect 16947 19068 17011 19072
rect 16947 19012 16951 19068
rect 16951 19012 17007 19068
rect 17007 19012 17011 19068
rect 16947 19008 17011 19012
rect 23009 19068 23073 19072
rect 23009 19012 23013 19068
rect 23013 19012 23069 19068
rect 23069 19012 23073 19068
rect 23009 19008 23073 19012
rect 23089 19068 23153 19072
rect 23089 19012 23093 19068
rect 23093 19012 23149 19068
rect 23149 19012 23153 19068
rect 23089 19008 23153 19012
rect 23169 19068 23233 19072
rect 23169 19012 23173 19068
rect 23173 19012 23229 19068
rect 23229 19012 23233 19068
rect 23169 19008 23233 19012
rect 23249 19068 23313 19072
rect 23249 19012 23253 19068
rect 23253 19012 23309 19068
rect 23309 19012 23313 19068
rect 23249 19008 23313 19012
rect 4763 18524 4827 18528
rect 4763 18468 4767 18524
rect 4767 18468 4823 18524
rect 4823 18468 4827 18524
rect 4763 18464 4827 18468
rect 4843 18524 4907 18528
rect 4843 18468 4847 18524
rect 4847 18468 4903 18524
rect 4903 18468 4907 18524
rect 4843 18464 4907 18468
rect 4923 18524 4987 18528
rect 4923 18468 4927 18524
rect 4927 18468 4983 18524
rect 4983 18468 4987 18524
rect 4923 18464 4987 18468
rect 5003 18524 5067 18528
rect 5003 18468 5007 18524
rect 5007 18468 5063 18524
rect 5063 18468 5067 18524
rect 5003 18464 5067 18468
rect 11065 18524 11129 18528
rect 11065 18468 11069 18524
rect 11069 18468 11125 18524
rect 11125 18468 11129 18524
rect 11065 18464 11129 18468
rect 11145 18524 11209 18528
rect 11145 18468 11149 18524
rect 11149 18468 11205 18524
rect 11205 18468 11209 18524
rect 11145 18464 11209 18468
rect 11225 18524 11289 18528
rect 11225 18468 11229 18524
rect 11229 18468 11285 18524
rect 11285 18468 11289 18524
rect 11225 18464 11289 18468
rect 11305 18524 11369 18528
rect 11305 18468 11309 18524
rect 11309 18468 11365 18524
rect 11365 18468 11369 18524
rect 11305 18464 11369 18468
rect 17367 18524 17431 18528
rect 17367 18468 17371 18524
rect 17371 18468 17427 18524
rect 17427 18468 17431 18524
rect 17367 18464 17431 18468
rect 17447 18524 17511 18528
rect 17447 18468 17451 18524
rect 17451 18468 17507 18524
rect 17507 18468 17511 18524
rect 17447 18464 17511 18468
rect 17527 18524 17591 18528
rect 17527 18468 17531 18524
rect 17531 18468 17587 18524
rect 17587 18468 17591 18524
rect 17527 18464 17591 18468
rect 17607 18524 17671 18528
rect 17607 18468 17611 18524
rect 17611 18468 17667 18524
rect 17667 18468 17671 18524
rect 17607 18464 17671 18468
rect 23669 18524 23733 18528
rect 23669 18468 23673 18524
rect 23673 18468 23729 18524
rect 23729 18468 23733 18524
rect 23669 18464 23733 18468
rect 23749 18524 23813 18528
rect 23749 18468 23753 18524
rect 23753 18468 23809 18524
rect 23809 18468 23813 18524
rect 23749 18464 23813 18468
rect 23829 18524 23893 18528
rect 23829 18468 23833 18524
rect 23833 18468 23889 18524
rect 23889 18468 23893 18524
rect 23829 18464 23893 18468
rect 23909 18524 23973 18528
rect 23909 18468 23913 18524
rect 23913 18468 23969 18524
rect 23969 18468 23973 18524
rect 23909 18464 23973 18468
rect 4103 17980 4167 17984
rect 4103 17924 4107 17980
rect 4107 17924 4163 17980
rect 4163 17924 4167 17980
rect 4103 17920 4167 17924
rect 4183 17980 4247 17984
rect 4183 17924 4187 17980
rect 4187 17924 4243 17980
rect 4243 17924 4247 17980
rect 4183 17920 4247 17924
rect 4263 17980 4327 17984
rect 4263 17924 4267 17980
rect 4267 17924 4323 17980
rect 4323 17924 4327 17980
rect 4263 17920 4327 17924
rect 4343 17980 4407 17984
rect 4343 17924 4347 17980
rect 4347 17924 4403 17980
rect 4403 17924 4407 17980
rect 4343 17920 4407 17924
rect 10405 17980 10469 17984
rect 10405 17924 10409 17980
rect 10409 17924 10465 17980
rect 10465 17924 10469 17980
rect 10405 17920 10469 17924
rect 10485 17980 10549 17984
rect 10485 17924 10489 17980
rect 10489 17924 10545 17980
rect 10545 17924 10549 17980
rect 10485 17920 10549 17924
rect 10565 17980 10629 17984
rect 10565 17924 10569 17980
rect 10569 17924 10625 17980
rect 10625 17924 10629 17980
rect 10565 17920 10629 17924
rect 10645 17980 10709 17984
rect 10645 17924 10649 17980
rect 10649 17924 10705 17980
rect 10705 17924 10709 17980
rect 10645 17920 10709 17924
rect 16707 17980 16771 17984
rect 16707 17924 16711 17980
rect 16711 17924 16767 17980
rect 16767 17924 16771 17980
rect 16707 17920 16771 17924
rect 16787 17980 16851 17984
rect 16787 17924 16791 17980
rect 16791 17924 16847 17980
rect 16847 17924 16851 17980
rect 16787 17920 16851 17924
rect 16867 17980 16931 17984
rect 16867 17924 16871 17980
rect 16871 17924 16927 17980
rect 16927 17924 16931 17980
rect 16867 17920 16931 17924
rect 16947 17980 17011 17984
rect 16947 17924 16951 17980
rect 16951 17924 17007 17980
rect 17007 17924 17011 17980
rect 16947 17920 17011 17924
rect 23009 17980 23073 17984
rect 23009 17924 23013 17980
rect 23013 17924 23069 17980
rect 23069 17924 23073 17980
rect 23009 17920 23073 17924
rect 23089 17980 23153 17984
rect 23089 17924 23093 17980
rect 23093 17924 23149 17980
rect 23149 17924 23153 17980
rect 23089 17920 23153 17924
rect 23169 17980 23233 17984
rect 23169 17924 23173 17980
rect 23173 17924 23229 17980
rect 23229 17924 23233 17980
rect 23169 17920 23233 17924
rect 23249 17980 23313 17984
rect 23249 17924 23253 17980
rect 23253 17924 23309 17980
rect 23309 17924 23313 17980
rect 23249 17920 23313 17924
rect 6132 17444 6196 17508
rect 4763 17436 4827 17440
rect 4763 17380 4767 17436
rect 4767 17380 4823 17436
rect 4823 17380 4827 17436
rect 4763 17376 4827 17380
rect 4843 17436 4907 17440
rect 4843 17380 4847 17436
rect 4847 17380 4903 17436
rect 4903 17380 4907 17436
rect 4843 17376 4907 17380
rect 4923 17436 4987 17440
rect 4923 17380 4927 17436
rect 4927 17380 4983 17436
rect 4983 17380 4987 17436
rect 4923 17376 4987 17380
rect 5003 17436 5067 17440
rect 5003 17380 5007 17436
rect 5007 17380 5063 17436
rect 5063 17380 5067 17436
rect 5003 17376 5067 17380
rect 11065 17436 11129 17440
rect 11065 17380 11069 17436
rect 11069 17380 11125 17436
rect 11125 17380 11129 17436
rect 11065 17376 11129 17380
rect 11145 17436 11209 17440
rect 11145 17380 11149 17436
rect 11149 17380 11205 17436
rect 11205 17380 11209 17436
rect 11145 17376 11209 17380
rect 11225 17436 11289 17440
rect 11225 17380 11229 17436
rect 11229 17380 11285 17436
rect 11285 17380 11289 17436
rect 11225 17376 11289 17380
rect 11305 17436 11369 17440
rect 11305 17380 11309 17436
rect 11309 17380 11365 17436
rect 11365 17380 11369 17436
rect 11305 17376 11369 17380
rect 17367 17436 17431 17440
rect 17367 17380 17371 17436
rect 17371 17380 17427 17436
rect 17427 17380 17431 17436
rect 17367 17376 17431 17380
rect 17447 17436 17511 17440
rect 17447 17380 17451 17436
rect 17451 17380 17507 17436
rect 17507 17380 17511 17436
rect 17447 17376 17511 17380
rect 17527 17436 17591 17440
rect 17527 17380 17531 17436
rect 17531 17380 17587 17436
rect 17587 17380 17591 17436
rect 17527 17376 17591 17380
rect 17607 17436 17671 17440
rect 17607 17380 17611 17436
rect 17611 17380 17667 17436
rect 17667 17380 17671 17436
rect 17607 17376 17671 17380
rect 23669 17436 23733 17440
rect 23669 17380 23673 17436
rect 23673 17380 23729 17436
rect 23729 17380 23733 17436
rect 23669 17376 23733 17380
rect 23749 17436 23813 17440
rect 23749 17380 23753 17436
rect 23753 17380 23809 17436
rect 23809 17380 23813 17436
rect 23749 17376 23813 17380
rect 23829 17436 23893 17440
rect 23829 17380 23833 17436
rect 23833 17380 23889 17436
rect 23889 17380 23893 17436
rect 23829 17376 23893 17380
rect 23909 17436 23973 17440
rect 23909 17380 23913 17436
rect 23913 17380 23969 17436
rect 23969 17380 23973 17436
rect 23909 17376 23973 17380
rect 4103 16892 4167 16896
rect 4103 16836 4107 16892
rect 4107 16836 4163 16892
rect 4163 16836 4167 16892
rect 4103 16832 4167 16836
rect 4183 16892 4247 16896
rect 4183 16836 4187 16892
rect 4187 16836 4243 16892
rect 4243 16836 4247 16892
rect 4183 16832 4247 16836
rect 4263 16892 4327 16896
rect 4263 16836 4267 16892
rect 4267 16836 4323 16892
rect 4323 16836 4327 16892
rect 4263 16832 4327 16836
rect 4343 16892 4407 16896
rect 4343 16836 4347 16892
rect 4347 16836 4403 16892
rect 4403 16836 4407 16892
rect 4343 16832 4407 16836
rect 10405 16892 10469 16896
rect 10405 16836 10409 16892
rect 10409 16836 10465 16892
rect 10465 16836 10469 16892
rect 10405 16832 10469 16836
rect 10485 16892 10549 16896
rect 10485 16836 10489 16892
rect 10489 16836 10545 16892
rect 10545 16836 10549 16892
rect 10485 16832 10549 16836
rect 10565 16892 10629 16896
rect 10565 16836 10569 16892
rect 10569 16836 10625 16892
rect 10625 16836 10629 16892
rect 10565 16832 10629 16836
rect 10645 16892 10709 16896
rect 10645 16836 10649 16892
rect 10649 16836 10705 16892
rect 10705 16836 10709 16892
rect 10645 16832 10709 16836
rect 16707 16892 16771 16896
rect 16707 16836 16711 16892
rect 16711 16836 16767 16892
rect 16767 16836 16771 16892
rect 16707 16832 16771 16836
rect 16787 16892 16851 16896
rect 16787 16836 16791 16892
rect 16791 16836 16847 16892
rect 16847 16836 16851 16892
rect 16787 16832 16851 16836
rect 16867 16892 16931 16896
rect 16867 16836 16871 16892
rect 16871 16836 16927 16892
rect 16927 16836 16931 16892
rect 16867 16832 16931 16836
rect 16947 16892 17011 16896
rect 16947 16836 16951 16892
rect 16951 16836 17007 16892
rect 17007 16836 17011 16892
rect 16947 16832 17011 16836
rect 23009 16892 23073 16896
rect 23009 16836 23013 16892
rect 23013 16836 23069 16892
rect 23069 16836 23073 16892
rect 23009 16832 23073 16836
rect 23089 16892 23153 16896
rect 23089 16836 23093 16892
rect 23093 16836 23149 16892
rect 23149 16836 23153 16892
rect 23089 16832 23153 16836
rect 23169 16892 23233 16896
rect 23169 16836 23173 16892
rect 23173 16836 23229 16892
rect 23229 16836 23233 16892
rect 23169 16832 23233 16836
rect 23249 16892 23313 16896
rect 23249 16836 23253 16892
rect 23253 16836 23309 16892
rect 23309 16836 23313 16892
rect 23249 16832 23313 16836
rect 4763 16348 4827 16352
rect 4763 16292 4767 16348
rect 4767 16292 4823 16348
rect 4823 16292 4827 16348
rect 4763 16288 4827 16292
rect 4843 16348 4907 16352
rect 4843 16292 4847 16348
rect 4847 16292 4903 16348
rect 4903 16292 4907 16348
rect 4843 16288 4907 16292
rect 4923 16348 4987 16352
rect 4923 16292 4927 16348
rect 4927 16292 4983 16348
rect 4983 16292 4987 16348
rect 4923 16288 4987 16292
rect 5003 16348 5067 16352
rect 5003 16292 5007 16348
rect 5007 16292 5063 16348
rect 5063 16292 5067 16348
rect 5003 16288 5067 16292
rect 11065 16348 11129 16352
rect 11065 16292 11069 16348
rect 11069 16292 11125 16348
rect 11125 16292 11129 16348
rect 11065 16288 11129 16292
rect 11145 16348 11209 16352
rect 11145 16292 11149 16348
rect 11149 16292 11205 16348
rect 11205 16292 11209 16348
rect 11145 16288 11209 16292
rect 11225 16348 11289 16352
rect 11225 16292 11229 16348
rect 11229 16292 11285 16348
rect 11285 16292 11289 16348
rect 11225 16288 11289 16292
rect 11305 16348 11369 16352
rect 11305 16292 11309 16348
rect 11309 16292 11365 16348
rect 11365 16292 11369 16348
rect 11305 16288 11369 16292
rect 17367 16348 17431 16352
rect 17367 16292 17371 16348
rect 17371 16292 17427 16348
rect 17427 16292 17431 16348
rect 17367 16288 17431 16292
rect 17447 16348 17511 16352
rect 17447 16292 17451 16348
rect 17451 16292 17507 16348
rect 17507 16292 17511 16348
rect 17447 16288 17511 16292
rect 17527 16348 17591 16352
rect 17527 16292 17531 16348
rect 17531 16292 17587 16348
rect 17587 16292 17591 16348
rect 17527 16288 17591 16292
rect 17607 16348 17671 16352
rect 17607 16292 17611 16348
rect 17611 16292 17667 16348
rect 17667 16292 17671 16348
rect 17607 16288 17671 16292
rect 23669 16348 23733 16352
rect 23669 16292 23673 16348
rect 23673 16292 23729 16348
rect 23729 16292 23733 16348
rect 23669 16288 23733 16292
rect 23749 16348 23813 16352
rect 23749 16292 23753 16348
rect 23753 16292 23809 16348
rect 23809 16292 23813 16348
rect 23749 16288 23813 16292
rect 23829 16348 23893 16352
rect 23829 16292 23833 16348
rect 23833 16292 23889 16348
rect 23889 16292 23893 16348
rect 23829 16288 23893 16292
rect 23909 16348 23973 16352
rect 23909 16292 23913 16348
rect 23913 16292 23969 16348
rect 23969 16292 23973 16348
rect 23909 16288 23973 16292
rect 4103 15804 4167 15808
rect 4103 15748 4107 15804
rect 4107 15748 4163 15804
rect 4163 15748 4167 15804
rect 4103 15744 4167 15748
rect 4183 15804 4247 15808
rect 4183 15748 4187 15804
rect 4187 15748 4243 15804
rect 4243 15748 4247 15804
rect 4183 15744 4247 15748
rect 4263 15804 4327 15808
rect 4263 15748 4267 15804
rect 4267 15748 4323 15804
rect 4323 15748 4327 15804
rect 4263 15744 4327 15748
rect 4343 15804 4407 15808
rect 4343 15748 4347 15804
rect 4347 15748 4403 15804
rect 4403 15748 4407 15804
rect 4343 15744 4407 15748
rect 10405 15804 10469 15808
rect 10405 15748 10409 15804
rect 10409 15748 10465 15804
rect 10465 15748 10469 15804
rect 10405 15744 10469 15748
rect 10485 15804 10549 15808
rect 10485 15748 10489 15804
rect 10489 15748 10545 15804
rect 10545 15748 10549 15804
rect 10485 15744 10549 15748
rect 10565 15804 10629 15808
rect 10565 15748 10569 15804
rect 10569 15748 10625 15804
rect 10625 15748 10629 15804
rect 10565 15744 10629 15748
rect 10645 15804 10709 15808
rect 10645 15748 10649 15804
rect 10649 15748 10705 15804
rect 10705 15748 10709 15804
rect 10645 15744 10709 15748
rect 16707 15804 16771 15808
rect 16707 15748 16711 15804
rect 16711 15748 16767 15804
rect 16767 15748 16771 15804
rect 16707 15744 16771 15748
rect 16787 15804 16851 15808
rect 16787 15748 16791 15804
rect 16791 15748 16847 15804
rect 16847 15748 16851 15804
rect 16787 15744 16851 15748
rect 16867 15804 16931 15808
rect 16867 15748 16871 15804
rect 16871 15748 16927 15804
rect 16927 15748 16931 15804
rect 16867 15744 16931 15748
rect 16947 15804 17011 15808
rect 16947 15748 16951 15804
rect 16951 15748 17007 15804
rect 17007 15748 17011 15804
rect 16947 15744 17011 15748
rect 23009 15804 23073 15808
rect 23009 15748 23013 15804
rect 23013 15748 23069 15804
rect 23069 15748 23073 15804
rect 23009 15744 23073 15748
rect 23089 15804 23153 15808
rect 23089 15748 23093 15804
rect 23093 15748 23149 15804
rect 23149 15748 23153 15804
rect 23089 15744 23153 15748
rect 23169 15804 23233 15808
rect 23169 15748 23173 15804
rect 23173 15748 23229 15804
rect 23229 15748 23233 15804
rect 23169 15744 23233 15748
rect 23249 15804 23313 15808
rect 23249 15748 23253 15804
rect 23253 15748 23309 15804
rect 23309 15748 23313 15804
rect 23249 15744 23313 15748
rect 4763 15260 4827 15264
rect 4763 15204 4767 15260
rect 4767 15204 4823 15260
rect 4823 15204 4827 15260
rect 4763 15200 4827 15204
rect 4843 15260 4907 15264
rect 4843 15204 4847 15260
rect 4847 15204 4903 15260
rect 4903 15204 4907 15260
rect 4843 15200 4907 15204
rect 4923 15260 4987 15264
rect 4923 15204 4927 15260
rect 4927 15204 4983 15260
rect 4983 15204 4987 15260
rect 4923 15200 4987 15204
rect 5003 15260 5067 15264
rect 5003 15204 5007 15260
rect 5007 15204 5063 15260
rect 5063 15204 5067 15260
rect 5003 15200 5067 15204
rect 11065 15260 11129 15264
rect 11065 15204 11069 15260
rect 11069 15204 11125 15260
rect 11125 15204 11129 15260
rect 11065 15200 11129 15204
rect 11145 15260 11209 15264
rect 11145 15204 11149 15260
rect 11149 15204 11205 15260
rect 11205 15204 11209 15260
rect 11145 15200 11209 15204
rect 11225 15260 11289 15264
rect 11225 15204 11229 15260
rect 11229 15204 11285 15260
rect 11285 15204 11289 15260
rect 11225 15200 11289 15204
rect 11305 15260 11369 15264
rect 11305 15204 11309 15260
rect 11309 15204 11365 15260
rect 11365 15204 11369 15260
rect 11305 15200 11369 15204
rect 17367 15260 17431 15264
rect 17367 15204 17371 15260
rect 17371 15204 17427 15260
rect 17427 15204 17431 15260
rect 17367 15200 17431 15204
rect 17447 15260 17511 15264
rect 17447 15204 17451 15260
rect 17451 15204 17507 15260
rect 17507 15204 17511 15260
rect 17447 15200 17511 15204
rect 17527 15260 17591 15264
rect 17527 15204 17531 15260
rect 17531 15204 17587 15260
rect 17587 15204 17591 15260
rect 17527 15200 17591 15204
rect 17607 15260 17671 15264
rect 17607 15204 17611 15260
rect 17611 15204 17667 15260
rect 17667 15204 17671 15260
rect 17607 15200 17671 15204
rect 23669 15260 23733 15264
rect 23669 15204 23673 15260
rect 23673 15204 23729 15260
rect 23729 15204 23733 15260
rect 23669 15200 23733 15204
rect 23749 15260 23813 15264
rect 23749 15204 23753 15260
rect 23753 15204 23809 15260
rect 23809 15204 23813 15260
rect 23749 15200 23813 15204
rect 23829 15260 23893 15264
rect 23829 15204 23833 15260
rect 23833 15204 23889 15260
rect 23889 15204 23893 15260
rect 23829 15200 23893 15204
rect 23909 15260 23973 15264
rect 23909 15204 23913 15260
rect 23913 15204 23969 15260
rect 23969 15204 23973 15260
rect 23909 15200 23973 15204
rect 5580 14996 5644 15060
rect 4103 14716 4167 14720
rect 4103 14660 4107 14716
rect 4107 14660 4163 14716
rect 4163 14660 4167 14716
rect 4103 14656 4167 14660
rect 4183 14716 4247 14720
rect 4183 14660 4187 14716
rect 4187 14660 4243 14716
rect 4243 14660 4247 14716
rect 4183 14656 4247 14660
rect 4263 14716 4327 14720
rect 4263 14660 4267 14716
rect 4267 14660 4323 14716
rect 4323 14660 4327 14716
rect 4263 14656 4327 14660
rect 4343 14716 4407 14720
rect 4343 14660 4347 14716
rect 4347 14660 4403 14716
rect 4403 14660 4407 14716
rect 4343 14656 4407 14660
rect 10405 14716 10469 14720
rect 10405 14660 10409 14716
rect 10409 14660 10465 14716
rect 10465 14660 10469 14716
rect 10405 14656 10469 14660
rect 10485 14716 10549 14720
rect 10485 14660 10489 14716
rect 10489 14660 10545 14716
rect 10545 14660 10549 14716
rect 10485 14656 10549 14660
rect 10565 14716 10629 14720
rect 10565 14660 10569 14716
rect 10569 14660 10625 14716
rect 10625 14660 10629 14716
rect 10565 14656 10629 14660
rect 10645 14716 10709 14720
rect 10645 14660 10649 14716
rect 10649 14660 10705 14716
rect 10705 14660 10709 14716
rect 10645 14656 10709 14660
rect 16707 14716 16771 14720
rect 16707 14660 16711 14716
rect 16711 14660 16767 14716
rect 16767 14660 16771 14716
rect 16707 14656 16771 14660
rect 16787 14716 16851 14720
rect 16787 14660 16791 14716
rect 16791 14660 16847 14716
rect 16847 14660 16851 14716
rect 16787 14656 16851 14660
rect 16867 14716 16931 14720
rect 16867 14660 16871 14716
rect 16871 14660 16927 14716
rect 16927 14660 16931 14716
rect 16867 14656 16931 14660
rect 16947 14716 17011 14720
rect 16947 14660 16951 14716
rect 16951 14660 17007 14716
rect 17007 14660 17011 14716
rect 16947 14656 17011 14660
rect 23009 14716 23073 14720
rect 23009 14660 23013 14716
rect 23013 14660 23069 14716
rect 23069 14660 23073 14716
rect 23009 14656 23073 14660
rect 23089 14716 23153 14720
rect 23089 14660 23093 14716
rect 23093 14660 23149 14716
rect 23149 14660 23153 14716
rect 23089 14656 23153 14660
rect 23169 14716 23233 14720
rect 23169 14660 23173 14716
rect 23173 14660 23229 14716
rect 23229 14660 23233 14716
rect 23169 14656 23233 14660
rect 23249 14716 23313 14720
rect 23249 14660 23253 14716
rect 23253 14660 23309 14716
rect 23309 14660 23313 14716
rect 23249 14656 23313 14660
rect 4763 14172 4827 14176
rect 4763 14116 4767 14172
rect 4767 14116 4823 14172
rect 4823 14116 4827 14172
rect 4763 14112 4827 14116
rect 4843 14172 4907 14176
rect 4843 14116 4847 14172
rect 4847 14116 4903 14172
rect 4903 14116 4907 14172
rect 4843 14112 4907 14116
rect 4923 14172 4987 14176
rect 4923 14116 4927 14172
rect 4927 14116 4983 14172
rect 4983 14116 4987 14172
rect 4923 14112 4987 14116
rect 5003 14172 5067 14176
rect 5003 14116 5007 14172
rect 5007 14116 5063 14172
rect 5063 14116 5067 14172
rect 5003 14112 5067 14116
rect 11065 14172 11129 14176
rect 11065 14116 11069 14172
rect 11069 14116 11125 14172
rect 11125 14116 11129 14172
rect 11065 14112 11129 14116
rect 11145 14172 11209 14176
rect 11145 14116 11149 14172
rect 11149 14116 11205 14172
rect 11205 14116 11209 14172
rect 11145 14112 11209 14116
rect 11225 14172 11289 14176
rect 11225 14116 11229 14172
rect 11229 14116 11285 14172
rect 11285 14116 11289 14172
rect 11225 14112 11289 14116
rect 11305 14172 11369 14176
rect 11305 14116 11309 14172
rect 11309 14116 11365 14172
rect 11365 14116 11369 14172
rect 11305 14112 11369 14116
rect 17367 14172 17431 14176
rect 17367 14116 17371 14172
rect 17371 14116 17427 14172
rect 17427 14116 17431 14172
rect 17367 14112 17431 14116
rect 17447 14172 17511 14176
rect 17447 14116 17451 14172
rect 17451 14116 17507 14172
rect 17507 14116 17511 14172
rect 17447 14112 17511 14116
rect 17527 14172 17591 14176
rect 17527 14116 17531 14172
rect 17531 14116 17587 14172
rect 17587 14116 17591 14172
rect 17527 14112 17591 14116
rect 17607 14172 17671 14176
rect 17607 14116 17611 14172
rect 17611 14116 17667 14172
rect 17667 14116 17671 14172
rect 17607 14112 17671 14116
rect 23669 14172 23733 14176
rect 23669 14116 23673 14172
rect 23673 14116 23729 14172
rect 23729 14116 23733 14172
rect 23669 14112 23733 14116
rect 23749 14172 23813 14176
rect 23749 14116 23753 14172
rect 23753 14116 23809 14172
rect 23809 14116 23813 14172
rect 23749 14112 23813 14116
rect 23829 14172 23893 14176
rect 23829 14116 23833 14172
rect 23833 14116 23889 14172
rect 23889 14116 23893 14172
rect 23829 14112 23893 14116
rect 23909 14172 23973 14176
rect 23909 14116 23913 14172
rect 23913 14116 23969 14172
rect 23969 14116 23973 14172
rect 23909 14112 23973 14116
rect 4103 13628 4167 13632
rect 4103 13572 4107 13628
rect 4107 13572 4163 13628
rect 4163 13572 4167 13628
rect 4103 13568 4167 13572
rect 4183 13628 4247 13632
rect 4183 13572 4187 13628
rect 4187 13572 4243 13628
rect 4243 13572 4247 13628
rect 4183 13568 4247 13572
rect 4263 13628 4327 13632
rect 4263 13572 4267 13628
rect 4267 13572 4323 13628
rect 4323 13572 4327 13628
rect 4263 13568 4327 13572
rect 4343 13628 4407 13632
rect 4343 13572 4347 13628
rect 4347 13572 4403 13628
rect 4403 13572 4407 13628
rect 4343 13568 4407 13572
rect 10405 13628 10469 13632
rect 10405 13572 10409 13628
rect 10409 13572 10465 13628
rect 10465 13572 10469 13628
rect 10405 13568 10469 13572
rect 10485 13628 10549 13632
rect 10485 13572 10489 13628
rect 10489 13572 10545 13628
rect 10545 13572 10549 13628
rect 10485 13568 10549 13572
rect 10565 13628 10629 13632
rect 10565 13572 10569 13628
rect 10569 13572 10625 13628
rect 10625 13572 10629 13628
rect 10565 13568 10629 13572
rect 10645 13628 10709 13632
rect 10645 13572 10649 13628
rect 10649 13572 10705 13628
rect 10705 13572 10709 13628
rect 10645 13568 10709 13572
rect 16707 13628 16771 13632
rect 16707 13572 16711 13628
rect 16711 13572 16767 13628
rect 16767 13572 16771 13628
rect 16707 13568 16771 13572
rect 16787 13628 16851 13632
rect 16787 13572 16791 13628
rect 16791 13572 16847 13628
rect 16847 13572 16851 13628
rect 16787 13568 16851 13572
rect 16867 13628 16931 13632
rect 16867 13572 16871 13628
rect 16871 13572 16927 13628
rect 16927 13572 16931 13628
rect 16867 13568 16931 13572
rect 16947 13628 17011 13632
rect 16947 13572 16951 13628
rect 16951 13572 17007 13628
rect 17007 13572 17011 13628
rect 16947 13568 17011 13572
rect 23009 13628 23073 13632
rect 23009 13572 23013 13628
rect 23013 13572 23069 13628
rect 23069 13572 23073 13628
rect 23009 13568 23073 13572
rect 23089 13628 23153 13632
rect 23089 13572 23093 13628
rect 23093 13572 23149 13628
rect 23149 13572 23153 13628
rect 23089 13568 23153 13572
rect 23169 13628 23233 13632
rect 23169 13572 23173 13628
rect 23173 13572 23229 13628
rect 23229 13572 23233 13628
rect 23169 13568 23233 13572
rect 23249 13628 23313 13632
rect 23249 13572 23253 13628
rect 23253 13572 23309 13628
rect 23309 13572 23313 13628
rect 23249 13568 23313 13572
rect 4763 13084 4827 13088
rect 4763 13028 4767 13084
rect 4767 13028 4823 13084
rect 4823 13028 4827 13084
rect 4763 13024 4827 13028
rect 4843 13084 4907 13088
rect 4843 13028 4847 13084
rect 4847 13028 4903 13084
rect 4903 13028 4907 13084
rect 4843 13024 4907 13028
rect 4923 13084 4987 13088
rect 4923 13028 4927 13084
rect 4927 13028 4983 13084
rect 4983 13028 4987 13084
rect 4923 13024 4987 13028
rect 5003 13084 5067 13088
rect 5003 13028 5007 13084
rect 5007 13028 5063 13084
rect 5063 13028 5067 13084
rect 5003 13024 5067 13028
rect 11065 13084 11129 13088
rect 11065 13028 11069 13084
rect 11069 13028 11125 13084
rect 11125 13028 11129 13084
rect 11065 13024 11129 13028
rect 11145 13084 11209 13088
rect 11145 13028 11149 13084
rect 11149 13028 11205 13084
rect 11205 13028 11209 13084
rect 11145 13024 11209 13028
rect 11225 13084 11289 13088
rect 11225 13028 11229 13084
rect 11229 13028 11285 13084
rect 11285 13028 11289 13084
rect 11225 13024 11289 13028
rect 11305 13084 11369 13088
rect 11305 13028 11309 13084
rect 11309 13028 11365 13084
rect 11365 13028 11369 13084
rect 11305 13024 11369 13028
rect 17367 13084 17431 13088
rect 17367 13028 17371 13084
rect 17371 13028 17427 13084
rect 17427 13028 17431 13084
rect 17367 13024 17431 13028
rect 17447 13084 17511 13088
rect 17447 13028 17451 13084
rect 17451 13028 17507 13084
rect 17507 13028 17511 13084
rect 17447 13024 17511 13028
rect 17527 13084 17591 13088
rect 17527 13028 17531 13084
rect 17531 13028 17587 13084
rect 17587 13028 17591 13084
rect 17527 13024 17591 13028
rect 17607 13084 17671 13088
rect 17607 13028 17611 13084
rect 17611 13028 17667 13084
rect 17667 13028 17671 13084
rect 17607 13024 17671 13028
rect 23669 13084 23733 13088
rect 23669 13028 23673 13084
rect 23673 13028 23729 13084
rect 23729 13028 23733 13084
rect 23669 13024 23733 13028
rect 23749 13084 23813 13088
rect 23749 13028 23753 13084
rect 23753 13028 23809 13084
rect 23809 13028 23813 13084
rect 23749 13024 23813 13028
rect 23829 13084 23893 13088
rect 23829 13028 23833 13084
rect 23833 13028 23889 13084
rect 23889 13028 23893 13084
rect 23829 13024 23893 13028
rect 23909 13084 23973 13088
rect 23909 13028 23913 13084
rect 23913 13028 23969 13084
rect 23969 13028 23973 13084
rect 23909 13024 23973 13028
rect 4103 12540 4167 12544
rect 4103 12484 4107 12540
rect 4107 12484 4163 12540
rect 4163 12484 4167 12540
rect 4103 12480 4167 12484
rect 4183 12540 4247 12544
rect 4183 12484 4187 12540
rect 4187 12484 4243 12540
rect 4243 12484 4247 12540
rect 4183 12480 4247 12484
rect 4263 12540 4327 12544
rect 4263 12484 4267 12540
rect 4267 12484 4323 12540
rect 4323 12484 4327 12540
rect 4263 12480 4327 12484
rect 4343 12540 4407 12544
rect 4343 12484 4347 12540
rect 4347 12484 4403 12540
rect 4403 12484 4407 12540
rect 4343 12480 4407 12484
rect 10405 12540 10469 12544
rect 10405 12484 10409 12540
rect 10409 12484 10465 12540
rect 10465 12484 10469 12540
rect 10405 12480 10469 12484
rect 10485 12540 10549 12544
rect 10485 12484 10489 12540
rect 10489 12484 10545 12540
rect 10545 12484 10549 12540
rect 10485 12480 10549 12484
rect 10565 12540 10629 12544
rect 10565 12484 10569 12540
rect 10569 12484 10625 12540
rect 10625 12484 10629 12540
rect 10565 12480 10629 12484
rect 10645 12540 10709 12544
rect 10645 12484 10649 12540
rect 10649 12484 10705 12540
rect 10705 12484 10709 12540
rect 10645 12480 10709 12484
rect 16707 12540 16771 12544
rect 16707 12484 16711 12540
rect 16711 12484 16767 12540
rect 16767 12484 16771 12540
rect 16707 12480 16771 12484
rect 16787 12540 16851 12544
rect 16787 12484 16791 12540
rect 16791 12484 16847 12540
rect 16847 12484 16851 12540
rect 16787 12480 16851 12484
rect 16867 12540 16931 12544
rect 16867 12484 16871 12540
rect 16871 12484 16927 12540
rect 16927 12484 16931 12540
rect 16867 12480 16931 12484
rect 16947 12540 17011 12544
rect 16947 12484 16951 12540
rect 16951 12484 17007 12540
rect 17007 12484 17011 12540
rect 16947 12480 17011 12484
rect 23009 12540 23073 12544
rect 23009 12484 23013 12540
rect 23013 12484 23069 12540
rect 23069 12484 23073 12540
rect 23009 12480 23073 12484
rect 23089 12540 23153 12544
rect 23089 12484 23093 12540
rect 23093 12484 23149 12540
rect 23149 12484 23153 12540
rect 23089 12480 23153 12484
rect 23169 12540 23233 12544
rect 23169 12484 23173 12540
rect 23173 12484 23229 12540
rect 23229 12484 23233 12540
rect 23169 12480 23233 12484
rect 23249 12540 23313 12544
rect 23249 12484 23253 12540
rect 23253 12484 23309 12540
rect 23309 12484 23313 12540
rect 23249 12480 23313 12484
rect 4763 11996 4827 12000
rect 4763 11940 4767 11996
rect 4767 11940 4823 11996
rect 4823 11940 4827 11996
rect 4763 11936 4827 11940
rect 4843 11996 4907 12000
rect 4843 11940 4847 11996
rect 4847 11940 4903 11996
rect 4903 11940 4907 11996
rect 4843 11936 4907 11940
rect 4923 11996 4987 12000
rect 4923 11940 4927 11996
rect 4927 11940 4983 11996
rect 4983 11940 4987 11996
rect 4923 11936 4987 11940
rect 5003 11996 5067 12000
rect 5003 11940 5007 11996
rect 5007 11940 5063 11996
rect 5063 11940 5067 11996
rect 5003 11936 5067 11940
rect 11065 11996 11129 12000
rect 11065 11940 11069 11996
rect 11069 11940 11125 11996
rect 11125 11940 11129 11996
rect 11065 11936 11129 11940
rect 11145 11996 11209 12000
rect 11145 11940 11149 11996
rect 11149 11940 11205 11996
rect 11205 11940 11209 11996
rect 11145 11936 11209 11940
rect 11225 11996 11289 12000
rect 11225 11940 11229 11996
rect 11229 11940 11285 11996
rect 11285 11940 11289 11996
rect 11225 11936 11289 11940
rect 11305 11996 11369 12000
rect 11305 11940 11309 11996
rect 11309 11940 11365 11996
rect 11365 11940 11369 11996
rect 11305 11936 11369 11940
rect 17367 11996 17431 12000
rect 17367 11940 17371 11996
rect 17371 11940 17427 11996
rect 17427 11940 17431 11996
rect 17367 11936 17431 11940
rect 17447 11996 17511 12000
rect 17447 11940 17451 11996
rect 17451 11940 17507 11996
rect 17507 11940 17511 11996
rect 17447 11936 17511 11940
rect 17527 11996 17591 12000
rect 17527 11940 17531 11996
rect 17531 11940 17587 11996
rect 17587 11940 17591 11996
rect 17527 11936 17591 11940
rect 17607 11996 17671 12000
rect 17607 11940 17611 11996
rect 17611 11940 17667 11996
rect 17667 11940 17671 11996
rect 17607 11936 17671 11940
rect 23669 11996 23733 12000
rect 23669 11940 23673 11996
rect 23673 11940 23729 11996
rect 23729 11940 23733 11996
rect 23669 11936 23733 11940
rect 23749 11996 23813 12000
rect 23749 11940 23753 11996
rect 23753 11940 23809 11996
rect 23809 11940 23813 11996
rect 23749 11936 23813 11940
rect 23829 11996 23893 12000
rect 23829 11940 23833 11996
rect 23833 11940 23889 11996
rect 23889 11940 23893 11996
rect 23829 11936 23893 11940
rect 23909 11996 23973 12000
rect 23909 11940 23913 11996
rect 23913 11940 23969 11996
rect 23969 11940 23973 11996
rect 23909 11936 23973 11940
rect 4103 11452 4167 11456
rect 4103 11396 4107 11452
rect 4107 11396 4163 11452
rect 4163 11396 4167 11452
rect 4103 11392 4167 11396
rect 4183 11452 4247 11456
rect 4183 11396 4187 11452
rect 4187 11396 4243 11452
rect 4243 11396 4247 11452
rect 4183 11392 4247 11396
rect 4263 11452 4327 11456
rect 4263 11396 4267 11452
rect 4267 11396 4323 11452
rect 4323 11396 4327 11452
rect 4263 11392 4327 11396
rect 4343 11452 4407 11456
rect 4343 11396 4347 11452
rect 4347 11396 4403 11452
rect 4403 11396 4407 11452
rect 4343 11392 4407 11396
rect 10405 11452 10469 11456
rect 10405 11396 10409 11452
rect 10409 11396 10465 11452
rect 10465 11396 10469 11452
rect 10405 11392 10469 11396
rect 10485 11452 10549 11456
rect 10485 11396 10489 11452
rect 10489 11396 10545 11452
rect 10545 11396 10549 11452
rect 10485 11392 10549 11396
rect 10565 11452 10629 11456
rect 10565 11396 10569 11452
rect 10569 11396 10625 11452
rect 10625 11396 10629 11452
rect 10565 11392 10629 11396
rect 10645 11452 10709 11456
rect 10645 11396 10649 11452
rect 10649 11396 10705 11452
rect 10705 11396 10709 11452
rect 10645 11392 10709 11396
rect 16707 11452 16771 11456
rect 16707 11396 16711 11452
rect 16711 11396 16767 11452
rect 16767 11396 16771 11452
rect 16707 11392 16771 11396
rect 16787 11452 16851 11456
rect 16787 11396 16791 11452
rect 16791 11396 16847 11452
rect 16847 11396 16851 11452
rect 16787 11392 16851 11396
rect 16867 11452 16931 11456
rect 16867 11396 16871 11452
rect 16871 11396 16927 11452
rect 16927 11396 16931 11452
rect 16867 11392 16931 11396
rect 16947 11452 17011 11456
rect 16947 11396 16951 11452
rect 16951 11396 17007 11452
rect 17007 11396 17011 11452
rect 16947 11392 17011 11396
rect 23009 11452 23073 11456
rect 23009 11396 23013 11452
rect 23013 11396 23069 11452
rect 23069 11396 23073 11452
rect 23009 11392 23073 11396
rect 23089 11452 23153 11456
rect 23089 11396 23093 11452
rect 23093 11396 23149 11452
rect 23149 11396 23153 11452
rect 23089 11392 23153 11396
rect 23169 11452 23233 11456
rect 23169 11396 23173 11452
rect 23173 11396 23229 11452
rect 23229 11396 23233 11452
rect 23169 11392 23233 11396
rect 23249 11452 23313 11456
rect 23249 11396 23253 11452
rect 23253 11396 23309 11452
rect 23309 11396 23313 11452
rect 23249 11392 23313 11396
rect 5580 11248 5644 11252
rect 5580 11192 5594 11248
rect 5594 11192 5644 11248
rect 5580 11188 5644 11192
rect 6316 11248 6380 11252
rect 6316 11192 6366 11248
rect 6366 11192 6380 11248
rect 6316 11188 6380 11192
rect 4763 10908 4827 10912
rect 4763 10852 4767 10908
rect 4767 10852 4823 10908
rect 4823 10852 4827 10908
rect 4763 10848 4827 10852
rect 4843 10908 4907 10912
rect 4843 10852 4847 10908
rect 4847 10852 4903 10908
rect 4903 10852 4907 10908
rect 4843 10848 4907 10852
rect 4923 10908 4987 10912
rect 4923 10852 4927 10908
rect 4927 10852 4983 10908
rect 4983 10852 4987 10908
rect 4923 10848 4987 10852
rect 5003 10908 5067 10912
rect 5003 10852 5007 10908
rect 5007 10852 5063 10908
rect 5063 10852 5067 10908
rect 5003 10848 5067 10852
rect 11065 10908 11129 10912
rect 11065 10852 11069 10908
rect 11069 10852 11125 10908
rect 11125 10852 11129 10908
rect 11065 10848 11129 10852
rect 11145 10908 11209 10912
rect 11145 10852 11149 10908
rect 11149 10852 11205 10908
rect 11205 10852 11209 10908
rect 11145 10848 11209 10852
rect 11225 10908 11289 10912
rect 11225 10852 11229 10908
rect 11229 10852 11285 10908
rect 11285 10852 11289 10908
rect 11225 10848 11289 10852
rect 11305 10908 11369 10912
rect 11305 10852 11309 10908
rect 11309 10852 11365 10908
rect 11365 10852 11369 10908
rect 11305 10848 11369 10852
rect 17367 10908 17431 10912
rect 17367 10852 17371 10908
rect 17371 10852 17427 10908
rect 17427 10852 17431 10908
rect 17367 10848 17431 10852
rect 17447 10908 17511 10912
rect 17447 10852 17451 10908
rect 17451 10852 17507 10908
rect 17507 10852 17511 10908
rect 17447 10848 17511 10852
rect 17527 10908 17591 10912
rect 17527 10852 17531 10908
rect 17531 10852 17587 10908
rect 17587 10852 17591 10908
rect 17527 10848 17591 10852
rect 17607 10908 17671 10912
rect 17607 10852 17611 10908
rect 17611 10852 17667 10908
rect 17667 10852 17671 10908
rect 17607 10848 17671 10852
rect 23669 10908 23733 10912
rect 23669 10852 23673 10908
rect 23673 10852 23729 10908
rect 23729 10852 23733 10908
rect 23669 10848 23733 10852
rect 23749 10908 23813 10912
rect 23749 10852 23753 10908
rect 23753 10852 23809 10908
rect 23809 10852 23813 10908
rect 23749 10848 23813 10852
rect 23829 10908 23893 10912
rect 23829 10852 23833 10908
rect 23833 10852 23889 10908
rect 23889 10852 23893 10908
rect 23829 10848 23893 10852
rect 23909 10908 23973 10912
rect 23909 10852 23913 10908
rect 23913 10852 23969 10908
rect 23969 10852 23973 10908
rect 23909 10848 23973 10852
rect 4103 10364 4167 10368
rect 4103 10308 4107 10364
rect 4107 10308 4163 10364
rect 4163 10308 4167 10364
rect 4103 10304 4167 10308
rect 4183 10364 4247 10368
rect 4183 10308 4187 10364
rect 4187 10308 4243 10364
rect 4243 10308 4247 10364
rect 4183 10304 4247 10308
rect 4263 10364 4327 10368
rect 4263 10308 4267 10364
rect 4267 10308 4323 10364
rect 4323 10308 4327 10364
rect 4263 10304 4327 10308
rect 4343 10364 4407 10368
rect 4343 10308 4347 10364
rect 4347 10308 4403 10364
rect 4403 10308 4407 10364
rect 4343 10304 4407 10308
rect 10405 10364 10469 10368
rect 10405 10308 10409 10364
rect 10409 10308 10465 10364
rect 10465 10308 10469 10364
rect 10405 10304 10469 10308
rect 10485 10364 10549 10368
rect 10485 10308 10489 10364
rect 10489 10308 10545 10364
rect 10545 10308 10549 10364
rect 10485 10304 10549 10308
rect 10565 10364 10629 10368
rect 10565 10308 10569 10364
rect 10569 10308 10625 10364
rect 10625 10308 10629 10364
rect 10565 10304 10629 10308
rect 10645 10364 10709 10368
rect 10645 10308 10649 10364
rect 10649 10308 10705 10364
rect 10705 10308 10709 10364
rect 10645 10304 10709 10308
rect 16707 10364 16771 10368
rect 16707 10308 16711 10364
rect 16711 10308 16767 10364
rect 16767 10308 16771 10364
rect 16707 10304 16771 10308
rect 16787 10364 16851 10368
rect 16787 10308 16791 10364
rect 16791 10308 16847 10364
rect 16847 10308 16851 10364
rect 16787 10304 16851 10308
rect 16867 10364 16931 10368
rect 16867 10308 16871 10364
rect 16871 10308 16927 10364
rect 16927 10308 16931 10364
rect 16867 10304 16931 10308
rect 16947 10364 17011 10368
rect 16947 10308 16951 10364
rect 16951 10308 17007 10364
rect 17007 10308 17011 10364
rect 16947 10304 17011 10308
rect 23009 10364 23073 10368
rect 23009 10308 23013 10364
rect 23013 10308 23069 10364
rect 23069 10308 23073 10364
rect 23009 10304 23073 10308
rect 23089 10364 23153 10368
rect 23089 10308 23093 10364
rect 23093 10308 23149 10364
rect 23149 10308 23153 10364
rect 23089 10304 23153 10308
rect 23169 10364 23233 10368
rect 23169 10308 23173 10364
rect 23173 10308 23229 10364
rect 23229 10308 23233 10364
rect 23169 10304 23233 10308
rect 23249 10364 23313 10368
rect 23249 10308 23253 10364
rect 23253 10308 23309 10364
rect 23309 10308 23313 10364
rect 23249 10304 23313 10308
rect 4763 9820 4827 9824
rect 4763 9764 4767 9820
rect 4767 9764 4823 9820
rect 4823 9764 4827 9820
rect 4763 9760 4827 9764
rect 4843 9820 4907 9824
rect 4843 9764 4847 9820
rect 4847 9764 4903 9820
rect 4903 9764 4907 9820
rect 4843 9760 4907 9764
rect 4923 9820 4987 9824
rect 4923 9764 4927 9820
rect 4927 9764 4983 9820
rect 4983 9764 4987 9820
rect 4923 9760 4987 9764
rect 5003 9820 5067 9824
rect 5003 9764 5007 9820
rect 5007 9764 5063 9820
rect 5063 9764 5067 9820
rect 5003 9760 5067 9764
rect 11065 9820 11129 9824
rect 11065 9764 11069 9820
rect 11069 9764 11125 9820
rect 11125 9764 11129 9820
rect 11065 9760 11129 9764
rect 11145 9820 11209 9824
rect 11145 9764 11149 9820
rect 11149 9764 11205 9820
rect 11205 9764 11209 9820
rect 11145 9760 11209 9764
rect 11225 9820 11289 9824
rect 11225 9764 11229 9820
rect 11229 9764 11285 9820
rect 11285 9764 11289 9820
rect 11225 9760 11289 9764
rect 11305 9820 11369 9824
rect 11305 9764 11309 9820
rect 11309 9764 11365 9820
rect 11365 9764 11369 9820
rect 11305 9760 11369 9764
rect 17367 9820 17431 9824
rect 17367 9764 17371 9820
rect 17371 9764 17427 9820
rect 17427 9764 17431 9820
rect 17367 9760 17431 9764
rect 17447 9820 17511 9824
rect 17447 9764 17451 9820
rect 17451 9764 17507 9820
rect 17507 9764 17511 9820
rect 17447 9760 17511 9764
rect 17527 9820 17591 9824
rect 17527 9764 17531 9820
rect 17531 9764 17587 9820
rect 17587 9764 17591 9820
rect 17527 9760 17591 9764
rect 17607 9820 17671 9824
rect 17607 9764 17611 9820
rect 17611 9764 17667 9820
rect 17667 9764 17671 9820
rect 17607 9760 17671 9764
rect 23669 9820 23733 9824
rect 23669 9764 23673 9820
rect 23673 9764 23729 9820
rect 23729 9764 23733 9820
rect 23669 9760 23733 9764
rect 23749 9820 23813 9824
rect 23749 9764 23753 9820
rect 23753 9764 23809 9820
rect 23809 9764 23813 9820
rect 23749 9760 23813 9764
rect 23829 9820 23893 9824
rect 23829 9764 23833 9820
rect 23833 9764 23889 9820
rect 23889 9764 23893 9820
rect 23829 9760 23893 9764
rect 23909 9820 23973 9824
rect 23909 9764 23913 9820
rect 23913 9764 23969 9820
rect 23969 9764 23973 9820
rect 23909 9760 23973 9764
rect 4103 9276 4167 9280
rect 4103 9220 4107 9276
rect 4107 9220 4163 9276
rect 4163 9220 4167 9276
rect 4103 9216 4167 9220
rect 4183 9276 4247 9280
rect 4183 9220 4187 9276
rect 4187 9220 4243 9276
rect 4243 9220 4247 9276
rect 4183 9216 4247 9220
rect 4263 9276 4327 9280
rect 4263 9220 4267 9276
rect 4267 9220 4323 9276
rect 4323 9220 4327 9276
rect 4263 9216 4327 9220
rect 4343 9276 4407 9280
rect 4343 9220 4347 9276
rect 4347 9220 4403 9276
rect 4403 9220 4407 9276
rect 4343 9216 4407 9220
rect 10405 9276 10469 9280
rect 10405 9220 10409 9276
rect 10409 9220 10465 9276
rect 10465 9220 10469 9276
rect 10405 9216 10469 9220
rect 10485 9276 10549 9280
rect 10485 9220 10489 9276
rect 10489 9220 10545 9276
rect 10545 9220 10549 9276
rect 10485 9216 10549 9220
rect 10565 9276 10629 9280
rect 10565 9220 10569 9276
rect 10569 9220 10625 9276
rect 10625 9220 10629 9276
rect 10565 9216 10629 9220
rect 10645 9276 10709 9280
rect 10645 9220 10649 9276
rect 10649 9220 10705 9276
rect 10705 9220 10709 9276
rect 10645 9216 10709 9220
rect 16707 9276 16771 9280
rect 16707 9220 16711 9276
rect 16711 9220 16767 9276
rect 16767 9220 16771 9276
rect 16707 9216 16771 9220
rect 16787 9276 16851 9280
rect 16787 9220 16791 9276
rect 16791 9220 16847 9276
rect 16847 9220 16851 9276
rect 16787 9216 16851 9220
rect 16867 9276 16931 9280
rect 16867 9220 16871 9276
rect 16871 9220 16927 9276
rect 16927 9220 16931 9276
rect 16867 9216 16931 9220
rect 16947 9276 17011 9280
rect 16947 9220 16951 9276
rect 16951 9220 17007 9276
rect 17007 9220 17011 9276
rect 16947 9216 17011 9220
rect 23009 9276 23073 9280
rect 23009 9220 23013 9276
rect 23013 9220 23069 9276
rect 23069 9220 23073 9276
rect 23009 9216 23073 9220
rect 23089 9276 23153 9280
rect 23089 9220 23093 9276
rect 23093 9220 23149 9276
rect 23149 9220 23153 9276
rect 23089 9216 23153 9220
rect 23169 9276 23233 9280
rect 23169 9220 23173 9276
rect 23173 9220 23229 9276
rect 23229 9220 23233 9276
rect 23169 9216 23233 9220
rect 23249 9276 23313 9280
rect 23249 9220 23253 9276
rect 23253 9220 23309 9276
rect 23309 9220 23313 9276
rect 23249 9216 23313 9220
rect 4763 8732 4827 8736
rect 4763 8676 4767 8732
rect 4767 8676 4823 8732
rect 4823 8676 4827 8732
rect 4763 8672 4827 8676
rect 4843 8732 4907 8736
rect 4843 8676 4847 8732
rect 4847 8676 4903 8732
rect 4903 8676 4907 8732
rect 4843 8672 4907 8676
rect 4923 8732 4987 8736
rect 4923 8676 4927 8732
rect 4927 8676 4983 8732
rect 4983 8676 4987 8732
rect 4923 8672 4987 8676
rect 5003 8732 5067 8736
rect 5003 8676 5007 8732
rect 5007 8676 5063 8732
rect 5063 8676 5067 8732
rect 5003 8672 5067 8676
rect 11065 8732 11129 8736
rect 11065 8676 11069 8732
rect 11069 8676 11125 8732
rect 11125 8676 11129 8732
rect 11065 8672 11129 8676
rect 11145 8732 11209 8736
rect 11145 8676 11149 8732
rect 11149 8676 11205 8732
rect 11205 8676 11209 8732
rect 11145 8672 11209 8676
rect 11225 8732 11289 8736
rect 11225 8676 11229 8732
rect 11229 8676 11285 8732
rect 11285 8676 11289 8732
rect 11225 8672 11289 8676
rect 11305 8732 11369 8736
rect 11305 8676 11309 8732
rect 11309 8676 11365 8732
rect 11365 8676 11369 8732
rect 11305 8672 11369 8676
rect 17367 8732 17431 8736
rect 17367 8676 17371 8732
rect 17371 8676 17427 8732
rect 17427 8676 17431 8732
rect 17367 8672 17431 8676
rect 17447 8732 17511 8736
rect 17447 8676 17451 8732
rect 17451 8676 17507 8732
rect 17507 8676 17511 8732
rect 17447 8672 17511 8676
rect 17527 8732 17591 8736
rect 17527 8676 17531 8732
rect 17531 8676 17587 8732
rect 17587 8676 17591 8732
rect 17527 8672 17591 8676
rect 17607 8732 17671 8736
rect 17607 8676 17611 8732
rect 17611 8676 17667 8732
rect 17667 8676 17671 8732
rect 17607 8672 17671 8676
rect 23669 8732 23733 8736
rect 23669 8676 23673 8732
rect 23673 8676 23729 8732
rect 23729 8676 23733 8732
rect 23669 8672 23733 8676
rect 23749 8732 23813 8736
rect 23749 8676 23753 8732
rect 23753 8676 23809 8732
rect 23809 8676 23813 8732
rect 23749 8672 23813 8676
rect 23829 8732 23893 8736
rect 23829 8676 23833 8732
rect 23833 8676 23889 8732
rect 23889 8676 23893 8732
rect 23829 8672 23893 8676
rect 23909 8732 23973 8736
rect 23909 8676 23913 8732
rect 23913 8676 23969 8732
rect 23969 8676 23973 8732
rect 23909 8672 23973 8676
rect 6316 8604 6380 8668
rect 4103 8188 4167 8192
rect 4103 8132 4107 8188
rect 4107 8132 4163 8188
rect 4163 8132 4167 8188
rect 4103 8128 4167 8132
rect 4183 8188 4247 8192
rect 4183 8132 4187 8188
rect 4187 8132 4243 8188
rect 4243 8132 4247 8188
rect 4183 8128 4247 8132
rect 4263 8188 4327 8192
rect 4263 8132 4267 8188
rect 4267 8132 4323 8188
rect 4323 8132 4327 8188
rect 4263 8128 4327 8132
rect 4343 8188 4407 8192
rect 4343 8132 4347 8188
rect 4347 8132 4403 8188
rect 4403 8132 4407 8188
rect 4343 8128 4407 8132
rect 10405 8188 10469 8192
rect 10405 8132 10409 8188
rect 10409 8132 10465 8188
rect 10465 8132 10469 8188
rect 10405 8128 10469 8132
rect 10485 8188 10549 8192
rect 10485 8132 10489 8188
rect 10489 8132 10545 8188
rect 10545 8132 10549 8188
rect 10485 8128 10549 8132
rect 10565 8188 10629 8192
rect 10565 8132 10569 8188
rect 10569 8132 10625 8188
rect 10625 8132 10629 8188
rect 10565 8128 10629 8132
rect 10645 8188 10709 8192
rect 10645 8132 10649 8188
rect 10649 8132 10705 8188
rect 10705 8132 10709 8188
rect 10645 8128 10709 8132
rect 16707 8188 16771 8192
rect 16707 8132 16711 8188
rect 16711 8132 16767 8188
rect 16767 8132 16771 8188
rect 16707 8128 16771 8132
rect 16787 8188 16851 8192
rect 16787 8132 16791 8188
rect 16791 8132 16847 8188
rect 16847 8132 16851 8188
rect 16787 8128 16851 8132
rect 16867 8188 16931 8192
rect 16867 8132 16871 8188
rect 16871 8132 16927 8188
rect 16927 8132 16931 8188
rect 16867 8128 16931 8132
rect 16947 8188 17011 8192
rect 16947 8132 16951 8188
rect 16951 8132 17007 8188
rect 17007 8132 17011 8188
rect 16947 8128 17011 8132
rect 23009 8188 23073 8192
rect 23009 8132 23013 8188
rect 23013 8132 23069 8188
rect 23069 8132 23073 8188
rect 23009 8128 23073 8132
rect 23089 8188 23153 8192
rect 23089 8132 23093 8188
rect 23093 8132 23149 8188
rect 23149 8132 23153 8188
rect 23089 8128 23153 8132
rect 23169 8188 23233 8192
rect 23169 8132 23173 8188
rect 23173 8132 23229 8188
rect 23229 8132 23233 8188
rect 23169 8128 23233 8132
rect 23249 8188 23313 8192
rect 23249 8132 23253 8188
rect 23253 8132 23309 8188
rect 23309 8132 23313 8188
rect 23249 8128 23313 8132
rect 5580 8120 5644 8124
rect 5580 8064 5630 8120
rect 5630 8064 5644 8120
rect 5580 8060 5644 8064
rect 4763 7644 4827 7648
rect 4763 7588 4767 7644
rect 4767 7588 4823 7644
rect 4823 7588 4827 7644
rect 4763 7584 4827 7588
rect 4843 7644 4907 7648
rect 4843 7588 4847 7644
rect 4847 7588 4903 7644
rect 4903 7588 4907 7644
rect 4843 7584 4907 7588
rect 4923 7644 4987 7648
rect 4923 7588 4927 7644
rect 4927 7588 4983 7644
rect 4983 7588 4987 7644
rect 4923 7584 4987 7588
rect 5003 7644 5067 7648
rect 5003 7588 5007 7644
rect 5007 7588 5063 7644
rect 5063 7588 5067 7644
rect 5003 7584 5067 7588
rect 11065 7644 11129 7648
rect 11065 7588 11069 7644
rect 11069 7588 11125 7644
rect 11125 7588 11129 7644
rect 11065 7584 11129 7588
rect 11145 7644 11209 7648
rect 11145 7588 11149 7644
rect 11149 7588 11205 7644
rect 11205 7588 11209 7644
rect 11145 7584 11209 7588
rect 11225 7644 11289 7648
rect 11225 7588 11229 7644
rect 11229 7588 11285 7644
rect 11285 7588 11289 7644
rect 11225 7584 11289 7588
rect 11305 7644 11369 7648
rect 11305 7588 11309 7644
rect 11309 7588 11365 7644
rect 11365 7588 11369 7644
rect 11305 7584 11369 7588
rect 17367 7644 17431 7648
rect 17367 7588 17371 7644
rect 17371 7588 17427 7644
rect 17427 7588 17431 7644
rect 17367 7584 17431 7588
rect 17447 7644 17511 7648
rect 17447 7588 17451 7644
rect 17451 7588 17507 7644
rect 17507 7588 17511 7644
rect 17447 7584 17511 7588
rect 17527 7644 17591 7648
rect 17527 7588 17531 7644
rect 17531 7588 17587 7644
rect 17587 7588 17591 7644
rect 17527 7584 17591 7588
rect 17607 7644 17671 7648
rect 17607 7588 17611 7644
rect 17611 7588 17667 7644
rect 17667 7588 17671 7644
rect 17607 7584 17671 7588
rect 23669 7644 23733 7648
rect 23669 7588 23673 7644
rect 23673 7588 23729 7644
rect 23729 7588 23733 7644
rect 23669 7584 23733 7588
rect 23749 7644 23813 7648
rect 23749 7588 23753 7644
rect 23753 7588 23809 7644
rect 23809 7588 23813 7644
rect 23749 7584 23813 7588
rect 23829 7644 23893 7648
rect 23829 7588 23833 7644
rect 23833 7588 23889 7644
rect 23889 7588 23893 7644
rect 23829 7584 23893 7588
rect 23909 7644 23973 7648
rect 23909 7588 23913 7644
rect 23913 7588 23969 7644
rect 23969 7588 23973 7644
rect 23909 7584 23973 7588
rect 4103 7100 4167 7104
rect 4103 7044 4107 7100
rect 4107 7044 4163 7100
rect 4163 7044 4167 7100
rect 4103 7040 4167 7044
rect 4183 7100 4247 7104
rect 4183 7044 4187 7100
rect 4187 7044 4243 7100
rect 4243 7044 4247 7100
rect 4183 7040 4247 7044
rect 4263 7100 4327 7104
rect 4263 7044 4267 7100
rect 4267 7044 4323 7100
rect 4323 7044 4327 7100
rect 4263 7040 4327 7044
rect 4343 7100 4407 7104
rect 4343 7044 4347 7100
rect 4347 7044 4403 7100
rect 4403 7044 4407 7100
rect 4343 7040 4407 7044
rect 10405 7100 10469 7104
rect 10405 7044 10409 7100
rect 10409 7044 10465 7100
rect 10465 7044 10469 7100
rect 10405 7040 10469 7044
rect 10485 7100 10549 7104
rect 10485 7044 10489 7100
rect 10489 7044 10545 7100
rect 10545 7044 10549 7100
rect 10485 7040 10549 7044
rect 10565 7100 10629 7104
rect 10565 7044 10569 7100
rect 10569 7044 10625 7100
rect 10625 7044 10629 7100
rect 10565 7040 10629 7044
rect 10645 7100 10709 7104
rect 10645 7044 10649 7100
rect 10649 7044 10705 7100
rect 10705 7044 10709 7100
rect 10645 7040 10709 7044
rect 16707 7100 16771 7104
rect 16707 7044 16711 7100
rect 16711 7044 16767 7100
rect 16767 7044 16771 7100
rect 16707 7040 16771 7044
rect 16787 7100 16851 7104
rect 16787 7044 16791 7100
rect 16791 7044 16847 7100
rect 16847 7044 16851 7100
rect 16787 7040 16851 7044
rect 16867 7100 16931 7104
rect 16867 7044 16871 7100
rect 16871 7044 16927 7100
rect 16927 7044 16931 7100
rect 16867 7040 16931 7044
rect 16947 7100 17011 7104
rect 16947 7044 16951 7100
rect 16951 7044 17007 7100
rect 17007 7044 17011 7100
rect 16947 7040 17011 7044
rect 23009 7100 23073 7104
rect 23009 7044 23013 7100
rect 23013 7044 23069 7100
rect 23069 7044 23073 7100
rect 23009 7040 23073 7044
rect 23089 7100 23153 7104
rect 23089 7044 23093 7100
rect 23093 7044 23149 7100
rect 23149 7044 23153 7100
rect 23089 7040 23153 7044
rect 23169 7100 23233 7104
rect 23169 7044 23173 7100
rect 23173 7044 23229 7100
rect 23229 7044 23233 7100
rect 23169 7040 23233 7044
rect 23249 7100 23313 7104
rect 23249 7044 23253 7100
rect 23253 7044 23309 7100
rect 23309 7044 23313 7100
rect 23249 7040 23313 7044
rect 4763 6556 4827 6560
rect 4763 6500 4767 6556
rect 4767 6500 4823 6556
rect 4823 6500 4827 6556
rect 4763 6496 4827 6500
rect 4843 6556 4907 6560
rect 4843 6500 4847 6556
rect 4847 6500 4903 6556
rect 4903 6500 4907 6556
rect 4843 6496 4907 6500
rect 4923 6556 4987 6560
rect 4923 6500 4927 6556
rect 4927 6500 4983 6556
rect 4983 6500 4987 6556
rect 4923 6496 4987 6500
rect 5003 6556 5067 6560
rect 5003 6500 5007 6556
rect 5007 6500 5063 6556
rect 5063 6500 5067 6556
rect 5003 6496 5067 6500
rect 11065 6556 11129 6560
rect 11065 6500 11069 6556
rect 11069 6500 11125 6556
rect 11125 6500 11129 6556
rect 11065 6496 11129 6500
rect 11145 6556 11209 6560
rect 11145 6500 11149 6556
rect 11149 6500 11205 6556
rect 11205 6500 11209 6556
rect 11145 6496 11209 6500
rect 11225 6556 11289 6560
rect 11225 6500 11229 6556
rect 11229 6500 11285 6556
rect 11285 6500 11289 6556
rect 11225 6496 11289 6500
rect 11305 6556 11369 6560
rect 11305 6500 11309 6556
rect 11309 6500 11365 6556
rect 11365 6500 11369 6556
rect 11305 6496 11369 6500
rect 17367 6556 17431 6560
rect 17367 6500 17371 6556
rect 17371 6500 17427 6556
rect 17427 6500 17431 6556
rect 17367 6496 17431 6500
rect 17447 6556 17511 6560
rect 17447 6500 17451 6556
rect 17451 6500 17507 6556
rect 17507 6500 17511 6556
rect 17447 6496 17511 6500
rect 17527 6556 17591 6560
rect 17527 6500 17531 6556
rect 17531 6500 17587 6556
rect 17587 6500 17591 6556
rect 17527 6496 17591 6500
rect 17607 6556 17671 6560
rect 17607 6500 17611 6556
rect 17611 6500 17667 6556
rect 17667 6500 17671 6556
rect 17607 6496 17671 6500
rect 23669 6556 23733 6560
rect 23669 6500 23673 6556
rect 23673 6500 23729 6556
rect 23729 6500 23733 6556
rect 23669 6496 23733 6500
rect 23749 6556 23813 6560
rect 23749 6500 23753 6556
rect 23753 6500 23809 6556
rect 23809 6500 23813 6556
rect 23749 6496 23813 6500
rect 23829 6556 23893 6560
rect 23829 6500 23833 6556
rect 23833 6500 23889 6556
rect 23889 6500 23893 6556
rect 23829 6496 23893 6500
rect 23909 6556 23973 6560
rect 23909 6500 23913 6556
rect 23913 6500 23969 6556
rect 23969 6500 23973 6556
rect 23909 6496 23973 6500
rect 4103 6012 4167 6016
rect 4103 5956 4107 6012
rect 4107 5956 4163 6012
rect 4163 5956 4167 6012
rect 4103 5952 4167 5956
rect 4183 6012 4247 6016
rect 4183 5956 4187 6012
rect 4187 5956 4243 6012
rect 4243 5956 4247 6012
rect 4183 5952 4247 5956
rect 4263 6012 4327 6016
rect 4263 5956 4267 6012
rect 4267 5956 4323 6012
rect 4323 5956 4327 6012
rect 4263 5952 4327 5956
rect 4343 6012 4407 6016
rect 4343 5956 4347 6012
rect 4347 5956 4403 6012
rect 4403 5956 4407 6012
rect 4343 5952 4407 5956
rect 10405 6012 10469 6016
rect 10405 5956 10409 6012
rect 10409 5956 10465 6012
rect 10465 5956 10469 6012
rect 10405 5952 10469 5956
rect 10485 6012 10549 6016
rect 10485 5956 10489 6012
rect 10489 5956 10545 6012
rect 10545 5956 10549 6012
rect 10485 5952 10549 5956
rect 10565 6012 10629 6016
rect 10565 5956 10569 6012
rect 10569 5956 10625 6012
rect 10625 5956 10629 6012
rect 10565 5952 10629 5956
rect 10645 6012 10709 6016
rect 10645 5956 10649 6012
rect 10649 5956 10705 6012
rect 10705 5956 10709 6012
rect 10645 5952 10709 5956
rect 16707 6012 16771 6016
rect 16707 5956 16711 6012
rect 16711 5956 16767 6012
rect 16767 5956 16771 6012
rect 16707 5952 16771 5956
rect 16787 6012 16851 6016
rect 16787 5956 16791 6012
rect 16791 5956 16847 6012
rect 16847 5956 16851 6012
rect 16787 5952 16851 5956
rect 16867 6012 16931 6016
rect 16867 5956 16871 6012
rect 16871 5956 16927 6012
rect 16927 5956 16931 6012
rect 16867 5952 16931 5956
rect 16947 6012 17011 6016
rect 16947 5956 16951 6012
rect 16951 5956 17007 6012
rect 17007 5956 17011 6012
rect 16947 5952 17011 5956
rect 23009 6012 23073 6016
rect 23009 5956 23013 6012
rect 23013 5956 23069 6012
rect 23069 5956 23073 6012
rect 23009 5952 23073 5956
rect 23089 6012 23153 6016
rect 23089 5956 23093 6012
rect 23093 5956 23149 6012
rect 23149 5956 23153 6012
rect 23089 5952 23153 5956
rect 23169 6012 23233 6016
rect 23169 5956 23173 6012
rect 23173 5956 23229 6012
rect 23229 5956 23233 6012
rect 23169 5952 23233 5956
rect 23249 6012 23313 6016
rect 23249 5956 23253 6012
rect 23253 5956 23309 6012
rect 23309 5956 23313 6012
rect 23249 5952 23313 5956
rect 4763 5468 4827 5472
rect 4763 5412 4767 5468
rect 4767 5412 4823 5468
rect 4823 5412 4827 5468
rect 4763 5408 4827 5412
rect 4843 5468 4907 5472
rect 4843 5412 4847 5468
rect 4847 5412 4903 5468
rect 4903 5412 4907 5468
rect 4843 5408 4907 5412
rect 4923 5468 4987 5472
rect 4923 5412 4927 5468
rect 4927 5412 4983 5468
rect 4983 5412 4987 5468
rect 4923 5408 4987 5412
rect 5003 5468 5067 5472
rect 5003 5412 5007 5468
rect 5007 5412 5063 5468
rect 5063 5412 5067 5468
rect 5003 5408 5067 5412
rect 11065 5468 11129 5472
rect 11065 5412 11069 5468
rect 11069 5412 11125 5468
rect 11125 5412 11129 5468
rect 11065 5408 11129 5412
rect 11145 5468 11209 5472
rect 11145 5412 11149 5468
rect 11149 5412 11205 5468
rect 11205 5412 11209 5468
rect 11145 5408 11209 5412
rect 11225 5468 11289 5472
rect 11225 5412 11229 5468
rect 11229 5412 11285 5468
rect 11285 5412 11289 5468
rect 11225 5408 11289 5412
rect 11305 5468 11369 5472
rect 11305 5412 11309 5468
rect 11309 5412 11365 5468
rect 11365 5412 11369 5468
rect 11305 5408 11369 5412
rect 17367 5468 17431 5472
rect 17367 5412 17371 5468
rect 17371 5412 17427 5468
rect 17427 5412 17431 5468
rect 17367 5408 17431 5412
rect 17447 5468 17511 5472
rect 17447 5412 17451 5468
rect 17451 5412 17507 5468
rect 17507 5412 17511 5468
rect 17447 5408 17511 5412
rect 17527 5468 17591 5472
rect 17527 5412 17531 5468
rect 17531 5412 17587 5468
rect 17587 5412 17591 5468
rect 17527 5408 17591 5412
rect 17607 5468 17671 5472
rect 17607 5412 17611 5468
rect 17611 5412 17667 5468
rect 17667 5412 17671 5468
rect 17607 5408 17671 5412
rect 23669 5468 23733 5472
rect 23669 5412 23673 5468
rect 23673 5412 23729 5468
rect 23729 5412 23733 5468
rect 23669 5408 23733 5412
rect 23749 5468 23813 5472
rect 23749 5412 23753 5468
rect 23753 5412 23809 5468
rect 23809 5412 23813 5468
rect 23749 5408 23813 5412
rect 23829 5468 23893 5472
rect 23829 5412 23833 5468
rect 23833 5412 23889 5468
rect 23889 5412 23893 5468
rect 23829 5408 23893 5412
rect 23909 5468 23973 5472
rect 23909 5412 23913 5468
rect 23913 5412 23969 5468
rect 23969 5412 23973 5468
rect 23909 5408 23973 5412
rect 4103 4924 4167 4928
rect 4103 4868 4107 4924
rect 4107 4868 4163 4924
rect 4163 4868 4167 4924
rect 4103 4864 4167 4868
rect 4183 4924 4247 4928
rect 4183 4868 4187 4924
rect 4187 4868 4243 4924
rect 4243 4868 4247 4924
rect 4183 4864 4247 4868
rect 4263 4924 4327 4928
rect 4263 4868 4267 4924
rect 4267 4868 4323 4924
rect 4323 4868 4327 4924
rect 4263 4864 4327 4868
rect 4343 4924 4407 4928
rect 4343 4868 4347 4924
rect 4347 4868 4403 4924
rect 4403 4868 4407 4924
rect 4343 4864 4407 4868
rect 10405 4924 10469 4928
rect 10405 4868 10409 4924
rect 10409 4868 10465 4924
rect 10465 4868 10469 4924
rect 10405 4864 10469 4868
rect 10485 4924 10549 4928
rect 10485 4868 10489 4924
rect 10489 4868 10545 4924
rect 10545 4868 10549 4924
rect 10485 4864 10549 4868
rect 10565 4924 10629 4928
rect 10565 4868 10569 4924
rect 10569 4868 10625 4924
rect 10625 4868 10629 4924
rect 10565 4864 10629 4868
rect 10645 4924 10709 4928
rect 10645 4868 10649 4924
rect 10649 4868 10705 4924
rect 10705 4868 10709 4924
rect 10645 4864 10709 4868
rect 16707 4924 16771 4928
rect 16707 4868 16711 4924
rect 16711 4868 16767 4924
rect 16767 4868 16771 4924
rect 16707 4864 16771 4868
rect 16787 4924 16851 4928
rect 16787 4868 16791 4924
rect 16791 4868 16847 4924
rect 16847 4868 16851 4924
rect 16787 4864 16851 4868
rect 16867 4924 16931 4928
rect 16867 4868 16871 4924
rect 16871 4868 16927 4924
rect 16927 4868 16931 4924
rect 16867 4864 16931 4868
rect 16947 4924 17011 4928
rect 16947 4868 16951 4924
rect 16951 4868 17007 4924
rect 17007 4868 17011 4924
rect 16947 4864 17011 4868
rect 23009 4924 23073 4928
rect 23009 4868 23013 4924
rect 23013 4868 23069 4924
rect 23069 4868 23073 4924
rect 23009 4864 23073 4868
rect 23089 4924 23153 4928
rect 23089 4868 23093 4924
rect 23093 4868 23149 4924
rect 23149 4868 23153 4924
rect 23089 4864 23153 4868
rect 23169 4924 23233 4928
rect 23169 4868 23173 4924
rect 23173 4868 23229 4924
rect 23229 4868 23233 4924
rect 23169 4864 23233 4868
rect 23249 4924 23313 4928
rect 23249 4868 23253 4924
rect 23253 4868 23309 4924
rect 23309 4868 23313 4924
rect 23249 4864 23313 4868
rect 4763 4380 4827 4384
rect 4763 4324 4767 4380
rect 4767 4324 4823 4380
rect 4823 4324 4827 4380
rect 4763 4320 4827 4324
rect 4843 4380 4907 4384
rect 4843 4324 4847 4380
rect 4847 4324 4903 4380
rect 4903 4324 4907 4380
rect 4843 4320 4907 4324
rect 4923 4380 4987 4384
rect 4923 4324 4927 4380
rect 4927 4324 4983 4380
rect 4983 4324 4987 4380
rect 4923 4320 4987 4324
rect 5003 4380 5067 4384
rect 5003 4324 5007 4380
rect 5007 4324 5063 4380
rect 5063 4324 5067 4380
rect 5003 4320 5067 4324
rect 11065 4380 11129 4384
rect 11065 4324 11069 4380
rect 11069 4324 11125 4380
rect 11125 4324 11129 4380
rect 11065 4320 11129 4324
rect 11145 4380 11209 4384
rect 11145 4324 11149 4380
rect 11149 4324 11205 4380
rect 11205 4324 11209 4380
rect 11145 4320 11209 4324
rect 11225 4380 11289 4384
rect 11225 4324 11229 4380
rect 11229 4324 11285 4380
rect 11285 4324 11289 4380
rect 11225 4320 11289 4324
rect 11305 4380 11369 4384
rect 11305 4324 11309 4380
rect 11309 4324 11365 4380
rect 11365 4324 11369 4380
rect 11305 4320 11369 4324
rect 17367 4380 17431 4384
rect 17367 4324 17371 4380
rect 17371 4324 17427 4380
rect 17427 4324 17431 4380
rect 17367 4320 17431 4324
rect 17447 4380 17511 4384
rect 17447 4324 17451 4380
rect 17451 4324 17507 4380
rect 17507 4324 17511 4380
rect 17447 4320 17511 4324
rect 17527 4380 17591 4384
rect 17527 4324 17531 4380
rect 17531 4324 17587 4380
rect 17587 4324 17591 4380
rect 17527 4320 17591 4324
rect 17607 4380 17671 4384
rect 17607 4324 17611 4380
rect 17611 4324 17667 4380
rect 17667 4324 17671 4380
rect 17607 4320 17671 4324
rect 23669 4380 23733 4384
rect 23669 4324 23673 4380
rect 23673 4324 23729 4380
rect 23729 4324 23733 4380
rect 23669 4320 23733 4324
rect 23749 4380 23813 4384
rect 23749 4324 23753 4380
rect 23753 4324 23809 4380
rect 23809 4324 23813 4380
rect 23749 4320 23813 4324
rect 23829 4380 23893 4384
rect 23829 4324 23833 4380
rect 23833 4324 23889 4380
rect 23889 4324 23893 4380
rect 23829 4320 23893 4324
rect 23909 4380 23973 4384
rect 23909 4324 23913 4380
rect 23913 4324 23969 4380
rect 23969 4324 23973 4380
rect 23909 4320 23973 4324
rect 4103 3836 4167 3840
rect 4103 3780 4107 3836
rect 4107 3780 4163 3836
rect 4163 3780 4167 3836
rect 4103 3776 4167 3780
rect 4183 3836 4247 3840
rect 4183 3780 4187 3836
rect 4187 3780 4243 3836
rect 4243 3780 4247 3836
rect 4183 3776 4247 3780
rect 4263 3836 4327 3840
rect 4263 3780 4267 3836
rect 4267 3780 4323 3836
rect 4323 3780 4327 3836
rect 4263 3776 4327 3780
rect 4343 3836 4407 3840
rect 4343 3780 4347 3836
rect 4347 3780 4403 3836
rect 4403 3780 4407 3836
rect 4343 3776 4407 3780
rect 10405 3836 10469 3840
rect 10405 3780 10409 3836
rect 10409 3780 10465 3836
rect 10465 3780 10469 3836
rect 10405 3776 10469 3780
rect 10485 3836 10549 3840
rect 10485 3780 10489 3836
rect 10489 3780 10545 3836
rect 10545 3780 10549 3836
rect 10485 3776 10549 3780
rect 10565 3836 10629 3840
rect 10565 3780 10569 3836
rect 10569 3780 10625 3836
rect 10625 3780 10629 3836
rect 10565 3776 10629 3780
rect 10645 3836 10709 3840
rect 10645 3780 10649 3836
rect 10649 3780 10705 3836
rect 10705 3780 10709 3836
rect 10645 3776 10709 3780
rect 16707 3836 16771 3840
rect 16707 3780 16711 3836
rect 16711 3780 16767 3836
rect 16767 3780 16771 3836
rect 16707 3776 16771 3780
rect 16787 3836 16851 3840
rect 16787 3780 16791 3836
rect 16791 3780 16847 3836
rect 16847 3780 16851 3836
rect 16787 3776 16851 3780
rect 16867 3836 16931 3840
rect 16867 3780 16871 3836
rect 16871 3780 16927 3836
rect 16927 3780 16931 3836
rect 16867 3776 16931 3780
rect 16947 3836 17011 3840
rect 16947 3780 16951 3836
rect 16951 3780 17007 3836
rect 17007 3780 17011 3836
rect 16947 3776 17011 3780
rect 23009 3836 23073 3840
rect 23009 3780 23013 3836
rect 23013 3780 23069 3836
rect 23069 3780 23073 3836
rect 23009 3776 23073 3780
rect 23089 3836 23153 3840
rect 23089 3780 23093 3836
rect 23093 3780 23149 3836
rect 23149 3780 23153 3836
rect 23089 3776 23153 3780
rect 23169 3836 23233 3840
rect 23169 3780 23173 3836
rect 23173 3780 23229 3836
rect 23229 3780 23233 3836
rect 23169 3776 23233 3780
rect 23249 3836 23313 3840
rect 23249 3780 23253 3836
rect 23253 3780 23309 3836
rect 23309 3780 23313 3836
rect 23249 3776 23313 3780
rect 4763 3292 4827 3296
rect 4763 3236 4767 3292
rect 4767 3236 4823 3292
rect 4823 3236 4827 3292
rect 4763 3232 4827 3236
rect 4843 3292 4907 3296
rect 4843 3236 4847 3292
rect 4847 3236 4903 3292
rect 4903 3236 4907 3292
rect 4843 3232 4907 3236
rect 4923 3292 4987 3296
rect 4923 3236 4927 3292
rect 4927 3236 4983 3292
rect 4983 3236 4987 3292
rect 4923 3232 4987 3236
rect 5003 3292 5067 3296
rect 5003 3236 5007 3292
rect 5007 3236 5063 3292
rect 5063 3236 5067 3292
rect 5003 3232 5067 3236
rect 11065 3292 11129 3296
rect 11065 3236 11069 3292
rect 11069 3236 11125 3292
rect 11125 3236 11129 3292
rect 11065 3232 11129 3236
rect 11145 3292 11209 3296
rect 11145 3236 11149 3292
rect 11149 3236 11205 3292
rect 11205 3236 11209 3292
rect 11145 3232 11209 3236
rect 11225 3292 11289 3296
rect 11225 3236 11229 3292
rect 11229 3236 11285 3292
rect 11285 3236 11289 3292
rect 11225 3232 11289 3236
rect 11305 3292 11369 3296
rect 11305 3236 11309 3292
rect 11309 3236 11365 3292
rect 11365 3236 11369 3292
rect 11305 3232 11369 3236
rect 17367 3292 17431 3296
rect 17367 3236 17371 3292
rect 17371 3236 17427 3292
rect 17427 3236 17431 3292
rect 17367 3232 17431 3236
rect 17447 3292 17511 3296
rect 17447 3236 17451 3292
rect 17451 3236 17507 3292
rect 17507 3236 17511 3292
rect 17447 3232 17511 3236
rect 17527 3292 17591 3296
rect 17527 3236 17531 3292
rect 17531 3236 17587 3292
rect 17587 3236 17591 3292
rect 17527 3232 17591 3236
rect 17607 3292 17671 3296
rect 17607 3236 17611 3292
rect 17611 3236 17667 3292
rect 17667 3236 17671 3292
rect 17607 3232 17671 3236
rect 23669 3292 23733 3296
rect 23669 3236 23673 3292
rect 23673 3236 23729 3292
rect 23729 3236 23733 3292
rect 23669 3232 23733 3236
rect 23749 3292 23813 3296
rect 23749 3236 23753 3292
rect 23753 3236 23809 3292
rect 23809 3236 23813 3292
rect 23749 3232 23813 3236
rect 23829 3292 23893 3296
rect 23829 3236 23833 3292
rect 23833 3236 23889 3292
rect 23889 3236 23893 3292
rect 23829 3232 23893 3236
rect 23909 3292 23973 3296
rect 23909 3236 23913 3292
rect 23913 3236 23969 3292
rect 23969 3236 23973 3292
rect 23909 3232 23973 3236
rect 4103 2748 4167 2752
rect 4103 2692 4107 2748
rect 4107 2692 4163 2748
rect 4163 2692 4167 2748
rect 4103 2688 4167 2692
rect 4183 2748 4247 2752
rect 4183 2692 4187 2748
rect 4187 2692 4243 2748
rect 4243 2692 4247 2748
rect 4183 2688 4247 2692
rect 4263 2748 4327 2752
rect 4263 2692 4267 2748
rect 4267 2692 4323 2748
rect 4323 2692 4327 2748
rect 4263 2688 4327 2692
rect 4343 2748 4407 2752
rect 4343 2692 4347 2748
rect 4347 2692 4403 2748
rect 4403 2692 4407 2748
rect 4343 2688 4407 2692
rect 10405 2748 10469 2752
rect 10405 2692 10409 2748
rect 10409 2692 10465 2748
rect 10465 2692 10469 2748
rect 10405 2688 10469 2692
rect 10485 2748 10549 2752
rect 10485 2692 10489 2748
rect 10489 2692 10545 2748
rect 10545 2692 10549 2748
rect 10485 2688 10549 2692
rect 10565 2748 10629 2752
rect 10565 2692 10569 2748
rect 10569 2692 10625 2748
rect 10625 2692 10629 2748
rect 10565 2688 10629 2692
rect 10645 2748 10709 2752
rect 10645 2692 10649 2748
rect 10649 2692 10705 2748
rect 10705 2692 10709 2748
rect 10645 2688 10709 2692
rect 16707 2748 16771 2752
rect 16707 2692 16711 2748
rect 16711 2692 16767 2748
rect 16767 2692 16771 2748
rect 16707 2688 16771 2692
rect 16787 2748 16851 2752
rect 16787 2692 16791 2748
rect 16791 2692 16847 2748
rect 16847 2692 16851 2748
rect 16787 2688 16851 2692
rect 16867 2748 16931 2752
rect 16867 2692 16871 2748
rect 16871 2692 16927 2748
rect 16927 2692 16931 2748
rect 16867 2688 16931 2692
rect 16947 2748 17011 2752
rect 16947 2692 16951 2748
rect 16951 2692 17007 2748
rect 17007 2692 17011 2748
rect 16947 2688 17011 2692
rect 23009 2748 23073 2752
rect 23009 2692 23013 2748
rect 23013 2692 23069 2748
rect 23069 2692 23073 2748
rect 23009 2688 23073 2692
rect 23089 2748 23153 2752
rect 23089 2692 23093 2748
rect 23093 2692 23149 2748
rect 23149 2692 23153 2748
rect 23089 2688 23153 2692
rect 23169 2748 23233 2752
rect 23169 2692 23173 2748
rect 23173 2692 23229 2748
rect 23229 2692 23233 2748
rect 23169 2688 23233 2692
rect 23249 2748 23313 2752
rect 23249 2692 23253 2748
rect 23253 2692 23309 2748
rect 23309 2692 23313 2748
rect 23249 2688 23313 2692
rect 4763 2204 4827 2208
rect 4763 2148 4767 2204
rect 4767 2148 4823 2204
rect 4823 2148 4827 2204
rect 4763 2144 4827 2148
rect 4843 2204 4907 2208
rect 4843 2148 4847 2204
rect 4847 2148 4903 2204
rect 4903 2148 4907 2204
rect 4843 2144 4907 2148
rect 4923 2204 4987 2208
rect 4923 2148 4927 2204
rect 4927 2148 4983 2204
rect 4983 2148 4987 2204
rect 4923 2144 4987 2148
rect 5003 2204 5067 2208
rect 5003 2148 5007 2204
rect 5007 2148 5063 2204
rect 5063 2148 5067 2204
rect 5003 2144 5067 2148
rect 11065 2204 11129 2208
rect 11065 2148 11069 2204
rect 11069 2148 11125 2204
rect 11125 2148 11129 2204
rect 11065 2144 11129 2148
rect 11145 2204 11209 2208
rect 11145 2148 11149 2204
rect 11149 2148 11205 2204
rect 11205 2148 11209 2204
rect 11145 2144 11209 2148
rect 11225 2204 11289 2208
rect 11225 2148 11229 2204
rect 11229 2148 11285 2204
rect 11285 2148 11289 2204
rect 11225 2144 11289 2148
rect 11305 2204 11369 2208
rect 11305 2148 11309 2204
rect 11309 2148 11365 2204
rect 11365 2148 11369 2204
rect 11305 2144 11369 2148
rect 17367 2204 17431 2208
rect 17367 2148 17371 2204
rect 17371 2148 17427 2204
rect 17427 2148 17431 2204
rect 17367 2144 17431 2148
rect 17447 2204 17511 2208
rect 17447 2148 17451 2204
rect 17451 2148 17507 2204
rect 17507 2148 17511 2204
rect 17447 2144 17511 2148
rect 17527 2204 17591 2208
rect 17527 2148 17531 2204
rect 17531 2148 17587 2204
rect 17587 2148 17591 2204
rect 17527 2144 17591 2148
rect 17607 2204 17671 2208
rect 17607 2148 17611 2204
rect 17611 2148 17667 2204
rect 17667 2148 17671 2204
rect 17607 2144 17671 2148
rect 23669 2204 23733 2208
rect 23669 2148 23673 2204
rect 23673 2148 23729 2204
rect 23729 2148 23733 2204
rect 23669 2144 23733 2148
rect 23749 2204 23813 2208
rect 23749 2148 23753 2204
rect 23753 2148 23809 2204
rect 23809 2148 23813 2204
rect 23749 2144 23813 2148
rect 23829 2204 23893 2208
rect 23829 2148 23833 2204
rect 23833 2148 23889 2204
rect 23889 2148 23893 2204
rect 23829 2144 23893 2148
rect 23909 2204 23973 2208
rect 23909 2148 23913 2204
rect 23913 2148 23969 2204
rect 23969 2148 23973 2204
rect 23909 2144 23973 2148
<< metal4 >>
rect 4095 26688 4415 27248
rect 4095 26624 4103 26688
rect 4167 26624 4183 26688
rect 4247 26624 4263 26688
rect 4327 26624 4343 26688
rect 4407 26624 4415 26688
rect 4095 25600 4415 26624
rect 4095 25536 4103 25600
rect 4167 25536 4183 25600
rect 4247 25536 4263 25600
rect 4327 25536 4343 25600
rect 4407 25536 4415 25600
rect 4095 24512 4415 25536
rect 4095 24448 4103 24512
rect 4167 24448 4183 24512
rect 4247 24448 4263 24512
rect 4327 24448 4343 24512
rect 4407 24448 4415 24512
rect 4095 24190 4415 24448
rect 4095 23954 4137 24190
rect 4373 23954 4415 24190
rect 4095 23424 4415 23954
rect 4095 23360 4103 23424
rect 4167 23360 4183 23424
rect 4247 23360 4263 23424
rect 4327 23360 4343 23424
rect 4407 23360 4415 23424
rect 4095 22336 4415 23360
rect 4095 22272 4103 22336
rect 4167 22272 4183 22336
rect 4247 22272 4263 22336
rect 4327 22272 4343 22336
rect 4407 22272 4415 22336
rect 4095 21248 4415 22272
rect 4095 21184 4103 21248
rect 4167 21184 4183 21248
rect 4247 21184 4263 21248
rect 4327 21184 4343 21248
rect 4407 21184 4415 21248
rect 4095 20160 4415 21184
rect 4095 20096 4103 20160
rect 4167 20096 4183 20160
rect 4247 20096 4263 20160
rect 4327 20096 4343 20160
rect 4407 20096 4415 20160
rect 4095 19072 4415 20096
rect 4095 19008 4103 19072
rect 4167 19008 4183 19072
rect 4247 19008 4263 19072
rect 4327 19008 4343 19072
rect 4407 19008 4415 19072
rect 4095 17984 4415 19008
rect 4095 17920 4103 17984
rect 4167 17934 4183 17984
rect 4247 17934 4263 17984
rect 4327 17934 4343 17984
rect 4407 17920 4415 17984
rect 4095 17698 4137 17920
rect 4373 17698 4415 17920
rect 4095 16896 4415 17698
rect 4095 16832 4103 16896
rect 4167 16832 4183 16896
rect 4247 16832 4263 16896
rect 4327 16832 4343 16896
rect 4407 16832 4415 16896
rect 4095 15808 4415 16832
rect 4095 15744 4103 15808
rect 4167 15744 4183 15808
rect 4247 15744 4263 15808
rect 4327 15744 4343 15808
rect 4407 15744 4415 15808
rect 4095 14720 4415 15744
rect 4095 14656 4103 14720
rect 4167 14656 4183 14720
rect 4247 14656 4263 14720
rect 4327 14656 4343 14720
rect 4407 14656 4415 14720
rect 4095 13632 4415 14656
rect 4095 13568 4103 13632
rect 4167 13568 4183 13632
rect 4247 13568 4263 13632
rect 4327 13568 4343 13632
rect 4407 13568 4415 13632
rect 4095 12544 4415 13568
rect 4095 12480 4103 12544
rect 4167 12480 4183 12544
rect 4247 12480 4263 12544
rect 4327 12480 4343 12544
rect 4407 12480 4415 12544
rect 4095 11678 4415 12480
rect 4095 11456 4137 11678
rect 4373 11456 4415 11678
rect 4095 11392 4103 11456
rect 4167 11392 4183 11442
rect 4247 11392 4263 11442
rect 4327 11392 4343 11442
rect 4407 11392 4415 11456
rect 4095 10368 4415 11392
rect 4095 10304 4103 10368
rect 4167 10304 4183 10368
rect 4247 10304 4263 10368
rect 4327 10304 4343 10368
rect 4407 10304 4415 10368
rect 4095 9280 4415 10304
rect 4095 9216 4103 9280
rect 4167 9216 4183 9280
rect 4247 9216 4263 9280
rect 4327 9216 4343 9280
rect 4407 9216 4415 9280
rect 4095 8192 4415 9216
rect 4095 8128 4103 8192
rect 4167 8128 4183 8192
rect 4247 8128 4263 8192
rect 4327 8128 4343 8192
rect 4407 8128 4415 8192
rect 4095 7104 4415 8128
rect 4095 7040 4103 7104
rect 4167 7040 4183 7104
rect 4247 7040 4263 7104
rect 4327 7040 4343 7104
rect 4407 7040 4415 7104
rect 4095 6016 4415 7040
rect 4095 5952 4103 6016
rect 4167 5952 4183 6016
rect 4247 5952 4263 6016
rect 4327 5952 4343 6016
rect 4407 5952 4415 6016
rect 4095 5422 4415 5952
rect 4095 5186 4137 5422
rect 4373 5186 4415 5422
rect 4095 4928 4415 5186
rect 4095 4864 4103 4928
rect 4167 4864 4183 4928
rect 4247 4864 4263 4928
rect 4327 4864 4343 4928
rect 4407 4864 4415 4928
rect 4095 3840 4415 4864
rect 4095 3776 4103 3840
rect 4167 3776 4183 3840
rect 4247 3776 4263 3840
rect 4327 3776 4343 3840
rect 4407 3776 4415 3840
rect 4095 2752 4415 3776
rect 4095 2688 4103 2752
rect 4167 2688 4183 2752
rect 4247 2688 4263 2752
rect 4327 2688 4343 2752
rect 4407 2688 4415 2752
rect 4095 2128 4415 2688
rect 4755 27232 5075 27248
rect 4755 27168 4763 27232
rect 4827 27168 4843 27232
rect 4907 27168 4923 27232
rect 4987 27168 5003 27232
rect 5067 27168 5075 27232
rect 4755 26144 5075 27168
rect 4755 26080 4763 26144
rect 4827 26080 4843 26144
rect 4907 26080 4923 26144
rect 4987 26080 5003 26144
rect 5067 26080 5075 26144
rect 4755 25056 5075 26080
rect 4755 24992 4763 25056
rect 4827 24992 4843 25056
rect 4907 24992 4923 25056
rect 4987 24992 5003 25056
rect 5067 24992 5075 25056
rect 4755 24850 5075 24992
rect 4755 24614 4797 24850
rect 5033 24614 5075 24850
rect 4755 23968 5075 24614
rect 4755 23904 4763 23968
rect 4827 23904 4843 23968
rect 4907 23904 4923 23968
rect 4987 23904 5003 23968
rect 5067 23904 5075 23968
rect 4755 22880 5075 23904
rect 10397 26688 10717 27248
rect 10397 26624 10405 26688
rect 10469 26624 10485 26688
rect 10549 26624 10565 26688
rect 10629 26624 10645 26688
rect 10709 26624 10717 26688
rect 10397 25600 10717 26624
rect 10397 25536 10405 25600
rect 10469 25536 10485 25600
rect 10549 25536 10565 25600
rect 10629 25536 10645 25600
rect 10709 25536 10717 25600
rect 10397 24512 10717 25536
rect 10397 24448 10405 24512
rect 10469 24448 10485 24512
rect 10549 24448 10565 24512
rect 10629 24448 10645 24512
rect 10709 24448 10717 24512
rect 10397 24190 10717 24448
rect 10397 23954 10439 24190
rect 10675 23954 10717 24190
rect 5579 23492 5645 23493
rect 5579 23428 5580 23492
rect 5644 23428 5645 23492
rect 5579 23427 5645 23428
rect 4755 22816 4763 22880
rect 4827 22816 4843 22880
rect 4907 22816 4923 22880
rect 4987 22816 5003 22880
rect 5067 22816 5075 22880
rect 4755 21792 5075 22816
rect 4755 21728 4763 21792
rect 4827 21728 4843 21792
rect 4907 21728 4923 21792
rect 4987 21728 5003 21792
rect 5067 21728 5075 21792
rect 4755 20704 5075 21728
rect 4755 20640 4763 20704
rect 4827 20640 4843 20704
rect 4907 20640 4923 20704
rect 4987 20640 5003 20704
rect 5067 20640 5075 20704
rect 4755 19616 5075 20640
rect 4755 19552 4763 19616
rect 4827 19552 4843 19616
rect 4907 19552 4923 19616
rect 4987 19552 5003 19616
rect 5067 19552 5075 19616
rect 4755 18594 5075 19552
rect 4755 18528 4797 18594
rect 5033 18528 5075 18594
rect 4755 18464 4763 18528
rect 5067 18464 5075 18528
rect 4755 18358 4797 18464
rect 5033 18358 5075 18464
rect 4755 17440 5075 18358
rect 4755 17376 4763 17440
rect 4827 17376 4843 17440
rect 4907 17376 4923 17440
rect 4987 17376 5003 17440
rect 5067 17376 5075 17440
rect 4755 16352 5075 17376
rect 4755 16288 4763 16352
rect 4827 16288 4843 16352
rect 4907 16288 4923 16352
rect 4987 16288 5003 16352
rect 5067 16288 5075 16352
rect 4755 15264 5075 16288
rect 4755 15200 4763 15264
rect 4827 15200 4843 15264
rect 4907 15200 4923 15264
rect 4987 15200 5003 15264
rect 5067 15200 5075 15264
rect 4755 14176 5075 15200
rect 5582 15061 5642 23427
rect 10397 23424 10717 23954
rect 10397 23360 10405 23424
rect 10469 23360 10485 23424
rect 10549 23360 10565 23424
rect 10629 23360 10645 23424
rect 10709 23360 10717 23424
rect 10397 22336 10717 23360
rect 10397 22272 10405 22336
rect 10469 22272 10485 22336
rect 10549 22272 10565 22336
rect 10629 22272 10645 22336
rect 10709 22272 10717 22336
rect 6131 21996 6197 21997
rect 6131 21932 6132 21996
rect 6196 21932 6197 21996
rect 6131 21931 6197 21932
rect 6134 17509 6194 21931
rect 10397 21248 10717 22272
rect 10397 21184 10405 21248
rect 10469 21184 10485 21248
rect 10549 21184 10565 21248
rect 10629 21184 10645 21248
rect 10709 21184 10717 21248
rect 10397 20160 10717 21184
rect 10397 20096 10405 20160
rect 10469 20096 10485 20160
rect 10549 20096 10565 20160
rect 10629 20096 10645 20160
rect 10709 20096 10717 20160
rect 10397 19072 10717 20096
rect 10397 19008 10405 19072
rect 10469 19008 10485 19072
rect 10549 19008 10565 19072
rect 10629 19008 10645 19072
rect 10709 19008 10717 19072
rect 10397 17984 10717 19008
rect 10397 17920 10405 17984
rect 10469 17934 10485 17984
rect 10549 17934 10565 17984
rect 10629 17934 10645 17984
rect 10709 17920 10717 17984
rect 10397 17698 10439 17920
rect 10675 17698 10717 17920
rect 6131 17508 6197 17509
rect 6131 17444 6132 17508
rect 6196 17444 6197 17508
rect 6131 17443 6197 17444
rect 10397 16896 10717 17698
rect 10397 16832 10405 16896
rect 10469 16832 10485 16896
rect 10549 16832 10565 16896
rect 10629 16832 10645 16896
rect 10709 16832 10717 16896
rect 10397 15808 10717 16832
rect 10397 15744 10405 15808
rect 10469 15744 10485 15808
rect 10549 15744 10565 15808
rect 10629 15744 10645 15808
rect 10709 15744 10717 15808
rect 5579 15060 5645 15061
rect 5579 14996 5580 15060
rect 5644 14996 5645 15060
rect 5579 14995 5645 14996
rect 4755 14112 4763 14176
rect 4827 14112 4843 14176
rect 4907 14112 4923 14176
rect 4987 14112 5003 14176
rect 5067 14112 5075 14176
rect 4755 13088 5075 14112
rect 4755 13024 4763 13088
rect 4827 13024 4843 13088
rect 4907 13024 4923 13088
rect 4987 13024 5003 13088
rect 5067 13024 5075 13088
rect 4755 12338 5075 13024
rect 4755 12102 4797 12338
rect 5033 12102 5075 12338
rect 4755 12000 5075 12102
rect 4755 11936 4763 12000
rect 4827 11936 4843 12000
rect 4907 11936 4923 12000
rect 4987 11936 5003 12000
rect 5067 11936 5075 12000
rect 4755 10912 5075 11936
rect 10397 14720 10717 15744
rect 10397 14656 10405 14720
rect 10469 14656 10485 14720
rect 10549 14656 10565 14720
rect 10629 14656 10645 14720
rect 10709 14656 10717 14720
rect 10397 13632 10717 14656
rect 10397 13568 10405 13632
rect 10469 13568 10485 13632
rect 10549 13568 10565 13632
rect 10629 13568 10645 13632
rect 10709 13568 10717 13632
rect 10397 12544 10717 13568
rect 10397 12480 10405 12544
rect 10469 12480 10485 12544
rect 10549 12480 10565 12544
rect 10629 12480 10645 12544
rect 10709 12480 10717 12544
rect 10397 11678 10717 12480
rect 10397 11456 10439 11678
rect 10675 11456 10717 11678
rect 10397 11392 10405 11456
rect 10469 11392 10485 11442
rect 10549 11392 10565 11442
rect 10629 11392 10645 11442
rect 10709 11392 10717 11456
rect 5579 11252 5645 11253
rect 5579 11188 5580 11252
rect 5644 11188 5645 11252
rect 5579 11187 5645 11188
rect 6315 11252 6381 11253
rect 6315 11188 6316 11252
rect 6380 11188 6381 11252
rect 6315 11187 6381 11188
rect 4755 10848 4763 10912
rect 4827 10848 4843 10912
rect 4907 10848 4923 10912
rect 4987 10848 5003 10912
rect 5067 10848 5075 10912
rect 4755 9824 5075 10848
rect 4755 9760 4763 9824
rect 4827 9760 4843 9824
rect 4907 9760 4923 9824
rect 4987 9760 5003 9824
rect 5067 9760 5075 9824
rect 4755 8736 5075 9760
rect 4755 8672 4763 8736
rect 4827 8672 4843 8736
rect 4907 8672 4923 8736
rect 4987 8672 5003 8736
rect 5067 8672 5075 8736
rect 4755 7648 5075 8672
rect 5582 8125 5642 11187
rect 6318 8669 6378 11187
rect 10397 10368 10717 11392
rect 10397 10304 10405 10368
rect 10469 10304 10485 10368
rect 10549 10304 10565 10368
rect 10629 10304 10645 10368
rect 10709 10304 10717 10368
rect 10397 9280 10717 10304
rect 10397 9216 10405 9280
rect 10469 9216 10485 9280
rect 10549 9216 10565 9280
rect 10629 9216 10645 9280
rect 10709 9216 10717 9280
rect 6315 8668 6381 8669
rect 6315 8604 6316 8668
rect 6380 8604 6381 8668
rect 6315 8603 6381 8604
rect 10397 8192 10717 9216
rect 10397 8128 10405 8192
rect 10469 8128 10485 8192
rect 10549 8128 10565 8192
rect 10629 8128 10645 8192
rect 10709 8128 10717 8192
rect 5579 8124 5645 8125
rect 5579 8060 5580 8124
rect 5644 8060 5645 8124
rect 5579 8059 5645 8060
rect 4755 7584 4763 7648
rect 4827 7584 4843 7648
rect 4907 7584 4923 7648
rect 4987 7584 5003 7648
rect 5067 7584 5075 7648
rect 4755 6560 5075 7584
rect 4755 6496 4763 6560
rect 4827 6496 4843 6560
rect 4907 6496 4923 6560
rect 4987 6496 5003 6560
rect 5067 6496 5075 6560
rect 4755 6082 5075 6496
rect 4755 5846 4797 6082
rect 5033 5846 5075 6082
rect 4755 5472 5075 5846
rect 4755 5408 4763 5472
rect 4827 5408 4843 5472
rect 4907 5408 4923 5472
rect 4987 5408 5003 5472
rect 5067 5408 5075 5472
rect 4755 4384 5075 5408
rect 4755 4320 4763 4384
rect 4827 4320 4843 4384
rect 4907 4320 4923 4384
rect 4987 4320 5003 4384
rect 5067 4320 5075 4384
rect 4755 3296 5075 4320
rect 4755 3232 4763 3296
rect 4827 3232 4843 3296
rect 4907 3232 4923 3296
rect 4987 3232 5003 3296
rect 5067 3232 5075 3296
rect 4755 2208 5075 3232
rect 4755 2144 4763 2208
rect 4827 2144 4843 2208
rect 4907 2144 4923 2208
rect 4987 2144 5003 2208
rect 5067 2144 5075 2208
rect 4755 2128 5075 2144
rect 10397 7104 10717 8128
rect 10397 7040 10405 7104
rect 10469 7040 10485 7104
rect 10549 7040 10565 7104
rect 10629 7040 10645 7104
rect 10709 7040 10717 7104
rect 10397 6016 10717 7040
rect 10397 5952 10405 6016
rect 10469 5952 10485 6016
rect 10549 5952 10565 6016
rect 10629 5952 10645 6016
rect 10709 5952 10717 6016
rect 10397 5422 10717 5952
rect 10397 5186 10439 5422
rect 10675 5186 10717 5422
rect 10397 4928 10717 5186
rect 10397 4864 10405 4928
rect 10469 4864 10485 4928
rect 10549 4864 10565 4928
rect 10629 4864 10645 4928
rect 10709 4864 10717 4928
rect 10397 3840 10717 4864
rect 10397 3776 10405 3840
rect 10469 3776 10485 3840
rect 10549 3776 10565 3840
rect 10629 3776 10645 3840
rect 10709 3776 10717 3840
rect 10397 2752 10717 3776
rect 10397 2688 10405 2752
rect 10469 2688 10485 2752
rect 10549 2688 10565 2752
rect 10629 2688 10645 2752
rect 10709 2688 10717 2752
rect 10397 2128 10717 2688
rect 11057 27232 11377 27248
rect 11057 27168 11065 27232
rect 11129 27168 11145 27232
rect 11209 27168 11225 27232
rect 11289 27168 11305 27232
rect 11369 27168 11377 27232
rect 11057 26144 11377 27168
rect 11057 26080 11065 26144
rect 11129 26080 11145 26144
rect 11209 26080 11225 26144
rect 11289 26080 11305 26144
rect 11369 26080 11377 26144
rect 11057 25056 11377 26080
rect 11057 24992 11065 25056
rect 11129 24992 11145 25056
rect 11209 24992 11225 25056
rect 11289 24992 11305 25056
rect 11369 24992 11377 25056
rect 11057 24850 11377 24992
rect 11057 24614 11099 24850
rect 11335 24614 11377 24850
rect 11057 23968 11377 24614
rect 11057 23904 11065 23968
rect 11129 23904 11145 23968
rect 11209 23904 11225 23968
rect 11289 23904 11305 23968
rect 11369 23904 11377 23968
rect 11057 22880 11377 23904
rect 11057 22816 11065 22880
rect 11129 22816 11145 22880
rect 11209 22816 11225 22880
rect 11289 22816 11305 22880
rect 11369 22816 11377 22880
rect 11057 21792 11377 22816
rect 11057 21728 11065 21792
rect 11129 21728 11145 21792
rect 11209 21728 11225 21792
rect 11289 21728 11305 21792
rect 11369 21728 11377 21792
rect 11057 20704 11377 21728
rect 11057 20640 11065 20704
rect 11129 20640 11145 20704
rect 11209 20640 11225 20704
rect 11289 20640 11305 20704
rect 11369 20640 11377 20704
rect 11057 19616 11377 20640
rect 11057 19552 11065 19616
rect 11129 19552 11145 19616
rect 11209 19552 11225 19616
rect 11289 19552 11305 19616
rect 11369 19552 11377 19616
rect 11057 18594 11377 19552
rect 11057 18528 11099 18594
rect 11335 18528 11377 18594
rect 11057 18464 11065 18528
rect 11369 18464 11377 18528
rect 11057 18358 11099 18464
rect 11335 18358 11377 18464
rect 11057 17440 11377 18358
rect 11057 17376 11065 17440
rect 11129 17376 11145 17440
rect 11209 17376 11225 17440
rect 11289 17376 11305 17440
rect 11369 17376 11377 17440
rect 11057 16352 11377 17376
rect 11057 16288 11065 16352
rect 11129 16288 11145 16352
rect 11209 16288 11225 16352
rect 11289 16288 11305 16352
rect 11369 16288 11377 16352
rect 11057 15264 11377 16288
rect 11057 15200 11065 15264
rect 11129 15200 11145 15264
rect 11209 15200 11225 15264
rect 11289 15200 11305 15264
rect 11369 15200 11377 15264
rect 11057 14176 11377 15200
rect 11057 14112 11065 14176
rect 11129 14112 11145 14176
rect 11209 14112 11225 14176
rect 11289 14112 11305 14176
rect 11369 14112 11377 14176
rect 11057 13088 11377 14112
rect 11057 13024 11065 13088
rect 11129 13024 11145 13088
rect 11209 13024 11225 13088
rect 11289 13024 11305 13088
rect 11369 13024 11377 13088
rect 11057 12338 11377 13024
rect 11057 12102 11099 12338
rect 11335 12102 11377 12338
rect 11057 12000 11377 12102
rect 11057 11936 11065 12000
rect 11129 11936 11145 12000
rect 11209 11936 11225 12000
rect 11289 11936 11305 12000
rect 11369 11936 11377 12000
rect 11057 10912 11377 11936
rect 11057 10848 11065 10912
rect 11129 10848 11145 10912
rect 11209 10848 11225 10912
rect 11289 10848 11305 10912
rect 11369 10848 11377 10912
rect 11057 9824 11377 10848
rect 11057 9760 11065 9824
rect 11129 9760 11145 9824
rect 11209 9760 11225 9824
rect 11289 9760 11305 9824
rect 11369 9760 11377 9824
rect 11057 8736 11377 9760
rect 11057 8672 11065 8736
rect 11129 8672 11145 8736
rect 11209 8672 11225 8736
rect 11289 8672 11305 8736
rect 11369 8672 11377 8736
rect 11057 7648 11377 8672
rect 11057 7584 11065 7648
rect 11129 7584 11145 7648
rect 11209 7584 11225 7648
rect 11289 7584 11305 7648
rect 11369 7584 11377 7648
rect 11057 6560 11377 7584
rect 11057 6496 11065 6560
rect 11129 6496 11145 6560
rect 11209 6496 11225 6560
rect 11289 6496 11305 6560
rect 11369 6496 11377 6560
rect 11057 6082 11377 6496
rect 11057 5846 11099 6082
rect 11335 5846 11377 6082
rect 11057 5472 11377 5846
rect 11057 5408 11065 5472
rect 11129 5408 11145 5472
rect 11209 5408 11225 5472
rect 11289 5408 11305 5472
rect 11369 5408 11377 5472
rect 11057 4384 11377 5408
rect 11057 4320 11065 4384
rect 11129 4320 11145 4384
rect 11209 4320 11225 4384
rect 11289 4320 11305 4384
rect 11369 4320 11377 4384
rect 11057 3296 11377 4320
rect 11057 3232 11065 3296
rect 11129 3232 11145 3296
rect 11209 3232 11225 3296
rect 11289 3232 11305 3296
rect 11369 3232 11377 3296
rect 11057 2208 11377 3232
rect 11057 2144 11065 2208
rect 11129 2144 11145 2208
rect 11209 2144 11225 2208
rect 11289 2144 11305 2208
rect 11369 2144 11377 2208
rect 11057 2128 11377 2144
rect 16699 26688 17019 27248
rect 16699 26624 16707 26688
rect 16771 26624 16787 26688
rect 16851 26624 16867 26688
rect 16931 26624 16947 26688
rect 17011 26624 17019 26688
rect 16699 25600 17019 26624
rect 16699 25536 16707 25600
rect 16771 25536 16787 25600
rect 16851 25536 16867 25600
rect 16931 25536 16947 25600
rect 17011 25536 17019 25600
rect 16699 24512 17019 25536
rect 16699 24448 16707 24512
rect 16771 24448 16787 24512
rect 16851 24448 16867 24512
rect 16931 24448 16947 24512
rect 17011 24448 17019 24512
rect 16699 24190 17019 24448
rect 16699 23954 16741 24190
rect 16977 23954 17019 24190
rect 16699 23424 17019 23954
rect 16699 23360 16707 23424
rect 16771 23360 16787 23424
rect 16851 23360 16867 23424
rect 16931 23360 16947 23424
rect 17011 23360 17019 23424
rect 16699 22336 17019 23360
rect 16699 22272 16707 22336
rect 16771 22272 16787 22336
rect 16851 22272 16867 22336
rect 16931 22272 16947 22336
rect 17011 22272 17019 22336
rect 16699 21248 17019 22272
rect 16699 21184 16707 21248
rect 16771 21184 16787 21248
rect 16851 21184 16867 21248
rect 16931 21184 16947 21248
rect 17011 21184 17019 21248
rect 16699 20160 17019 21184
rect 16699 20096 16707 20160
rect 16771 20096 16787 20160
rect 16851 20096 16867 20160
rect 16931 20096 16947 20160
rect 17011 20096 17019 20160
rect 16699 19072 17019 20096
rect 16699 19008 16707 19072
rect 16771 19008 16787 19072
rect 16851 19008 16867 19072
rect 16931 19008 16947 19072
rect 17011 19008 17019 19072
rect 16699 17984 17019 19008
rect 16699 17920 16707 17984
rect 16771 17934 16787 17984
rect 16851 17934 16867 17984
rect 16931 17934 16947 17984
rect 17011 17920 17019 17984
rect 16699 17698 16741 17920
rect 16977 17698 17019 17920
rect 16699 16896 17019 17698
rect 16699 16832 16707 16896
rect 16771 16832 16787 16896
rect 16851 16832 16867 16896
rect 16931 16832 16947 16896
rect 17011 16832 17019 16896
rect 16699 15808 17019 16832
rect 16699 15744 16707 15808
rect 16771 15744 16787 15808
rect 16851 15744 16867 15808
rect 16931 15744 16947 15808
rect 17011 15744 17019 15808
rect 16699 14720 17019 15744
rect 16699 14656 16707 14720
rect 16771 14656 16787 14720
rect 16851 14656 16867 14720
rect 16931 14656 16947 14720
rect 17011 14656 17019 14720
rect 16699 13632 17019 14656
rect 16699 13568 16707 13632
rect 16771 13568 16787 13632
rect 16851 13568 16867 13632
rect 16931 13568 16947 13632
rect 17011 13568 17019 13632
rect 16699 12544 17019 13568
rect 16699 12480 16707 12544
rect 16771 12480 16787 12544
rect 16851 12480 16867 12544
rect 16931 12480 16947 12544
rect 17011 12480 17019 12544
rect 16699 11678 17019 12480
rect 16699 11456 16741 11678
rect 16977 11456 17019 11678
rect 16699 11392 16707 11456
rect 16771 11392 16787 11442
rect 16851 11392 16867 11442
rect 16931 11392 16947 11442
rect 17011 11392 17019 11456
rect 16699 10368 17019 11392
rect 16699 10304 16707 10368
rect 16771 10304 16787 10368
rect 16851 10304 16867 10368
rect 16931 10304 16947 10368
rect 17011 10304 17019 10368
rect 16699 9280 17019 10304
rect 16699 9216 16707 9280
rect 16771 9216 16787 9280
rect 16851 9216 16867 9280
rect 16931 9216 16947 9280
rect 17011 9216 17019 9280
rect 16699 8192 17019 9216
rect 16699 8128 16707 8192
rect 16771 8128 16787 8192
rect 16851 8128 16867 8192
rect 16931 8128 16947 8192
rect 17011 8128 17019 8192
rect 16699 7104 17019 8128
rect 16699 7040 16707 7104
rect 16771 7040 16787 7104
rect 16851 7040 16867 7104
rect 16931 7040 16947 7104
rect 17011 7040 17019 7104
rect 16699 6016 17019 7040
rect 16699 5952 16707 6016
rect 16771 5952 16787 6016
rect 16851 5952 16867 6016
rect 16931 5952 16947 6016
rect 17011 5952 17019 6016
rect 16699 5422 17019 5952
rect 16699 5186 16741 5422
rect 16977 5186 17019 5422
rect 16699 4928 17019 5186
rect 16699 4864 16707 4928
rect 16771 4864 16787 4928
rect 16851 4864 16867 4928
rect 16931 4864 16947 4928
rect 17011 4864 17019 4928
rect 16699 3840 17019 4864
rect 16699 3776 16707 3840
rect 16771 3776 16787 3840
rect 16851 3776 16867 3840
rect 16931 3776 16947 3840
rect 17011 3776 17019 3840
rect 16699 2752 17019 3776
rect 16699 2688 16707 2752
rect 16771 2688 16787 2752
rect 16851 2688 16867 2752
rect 16931 2688 16947 2752
rect 17011 2688 17019 2752
rect 16699 2128 17019 2688
rect 17359 27232 17679 27248
rect 17359 27168 17367 27232
rect 17431 27168 17447 27232
rect 17511 27168 17527 27232
rect 17591 27168 17607 27232
rect 17671 27168 17679 27232
rect 17359 26144 17679 27168
rect 17359 26080 17367 26144
rect 17431 26080 17447 26144
rect 17511 26080 17527 26144
rect 17591 26080 17607 26144
rect 17671 26080 17679 26144
rect 17359 25056 17679 26080
rect 17359 24992 17367 25056
rect 17431 24992 17447 25056
rect 17511 24992 17527 25056
rect 17591 24992 17607 25056
rect 17671 24992 17679 25056
rect 17359 24850 17679 24992
rect 17359 24614 17401 24850
rect 17637 24614 17679 24850
rect 17359 23968 17679 24614
rect 17359 23904 17367 23968
rect 17431 23904 17447 23968
rect 17511 23904 17527 23968
rect 17591 23904 17607 23968
rect 17671 23904 17679 23968
rect 17359 22880 17679 23904
rect 17359 22816 17367 22880
rect 17431 22816 17447 22880
rect 17511 22816 17527 22880
rect 17591 22816 17607 22880
rect 17671 22816 17679 22880
rect 17359 21792 17679 22816
rect 17359 21728 17367 21792
rect 17431 21728 17447 21792
rect 17511 21728 17527 21792
rect 17591 21728 17607 21792
rect 17671 21728 17679 21792
rect 17359 20704 17679 21728
rect 17359 20640 17367 20704
rect 17431 20640 17447 20704
rect 17511 20640 17527 20704
rect 17591 20640 17607 20704
rect 17671 20640 17679 20704
rect 17359 19616 17679 20640
rect 17359 19552 17367 19616
rect 17431 19552 17447 19616
rect 17511 19552 17527 19616
rect 17591 19552 17607 19616
rect 17671 19552 17679 19616
rect 17359 18594 17679 19552
rect 17359 18528 17401 18594
rect 17637 18528 17679 18594
rect 17359 18464 17367 18528
rect 17671 18464 17679 18528
rect 17359 18358 17401 18464
rect 17637 18358 17679 18464
rect 17359 17440 17679 18358
rect 17359 17376 17367 17440
rect 17431 17376 17447 17440
rect 17511 17376 17527 17440
rect 17591 17376 17607 17440
rect 17671 17376 17679 17440
rect 17359 16352 17679 17376
rect 17359 16288 17367 16352
rect 17431 16288 17447 16352
rect 17511 16288 17527 16352
rect 17591 16288 17607 16352
rect 17671 16288 17679 16352
rect 17359 15264 17679 16288
rect 17359 15200 17367 15264
rect 17431 15200 17447 15264
rect 17511 15200 17527 15264
rect 17591 15200 17607 15264
rect 17671 15200 17679 15264
rect 17359 14176 17679 15200
rect 17359 14112 17367 14176
rect 17431 14112 17447 14176
rect 17511 14112 17527 14176
rect 17591 14112 17607 14176
rect 17671 14112 17679 14176
rect 17359 13088 17679 14112
rect 17359 13024 17367 13088
rect 17431 13024 17447 13088
rect 17511 13024 17527 13088
rect 17591 13024 17607 13088
rect 17671 13024 17679 13088
rect 17359 12338 17679 13024
rect 17359 12102 17401 12338
rect 17637 12102 17679 12338
rect 17359 12000 17679 12102
rect 17359 11936 17367 12000
rect 17431 11936 17447 12000
rect 17511 11936 17527 12000
rect 17591 11936 17607 12000
rect 17671 11936 17679 12000
rect 17359 10912 17679 11936
rect 17359 10848 17367 10912
rect 17431 10848 17447 10912
rect 17511 10848 17527 10912
rect 17591 10848 17607 10912
rect 17671 10848 17679 10912
rect 17359 9824 17679 10848
rect 17359 9760 17367 9824
rect 17431 9760 17447 9824
rect 17511 9760 17527 9824
rect 17591 9760 17607 9824
rect 17671 9760 17679 9824
rect 17359 8736 17679 9760
rect 17359 8672 17367 8736
rect 17431 8672 17447 8736
rect 17511 8672 17527 8736
rect 17591 8672 17607 8736
rect 17671 8672 17679 8736
rect 17359 7648 17679 8672
rect 17359 7584 17367 7648
rect 17431 7584 17447 7648
rect 17511 7584 17527 7648
rect 17591 7584 17607 7648
rect 17671 7584 17679 7648
rect 17359 6560 17679 7584
rect 17359 6496 17367 6560
rect 17431 6496 17447 6560
rect 17511 6496 17527 6560
rect 17591 6496 17607 6560
rect 17671 6496 17679 6560
rect 17359 6082 17679 6496
rect 17359 5846 17401 6082
rect 17637 5846 17679 6082
rect 17359 5472 17679 5846
rect 17359 5408 17367 5472
rect 17431 5408 17447 5472
rect 17511 5408 17527 5472
rect 17591 5408 17607 5472
rect 17671 5408 17679 5472
rect 17359 4384 17679 5408
rect 17359 4320 17367 4384
rect 17431 4320 17447 4384
rect 17511 4320 17527 4384
rect 17591 4320 17607 4384
rect 17671 4320 17679 4384
rect 17359 3296 17679 4320
rect 17359 3232 17367 3296
rect 17431 3232 17447 3296
rect 17511 3232 17527 3296
rect 17591 3232 17607 3296
rect 17671 3232 17679 3296
rect 17359 2208 17679 3232
rect 17359 2144 17367 2208
rect 17431 2144 17447 2208
rect 17511 2144 17527 2208
rect 17591 2144 17607 2208
rect 17671 2144 17679 2208
rect 17359 2128 17679 2144
rect 23001 26688 23321 27248
rect 23001 26624 23009 26688
rect 23073 26624 23089 26688
rect 23153 26624 23169 26688
rect 23233 26624 23249 26688
rect 23313 26624 23321 26688
rect 23001 25600 23321 26624
rect 23001 25536 23009 25600
rect 23073 25536 23089 25600
rect 23153 25536 23169 25600
rect 23233 25536 23249 25600
rect 23313 25536 23321 25600
rect 23001 24512 23321 25536
rect 23001 24448 23009 24512
rect 23073 24448 23089 24512
rect 23153 24448 23169 24512
rect 23233 24448 23249 24512
rect 23313 24448 23321 24512
rect 23001 24190 23321 24448
rect 23001 23954 23043 24190
rect 23279 23954 23321 24190
rect 23001 23424 23321 23954
rect 23001 23360 23009 23424
rect 23073 23360 23089 23424
rect 23153 23360 23169 23424
rect 23233 23360 23249 23424
rect 23313 23360 23321 23424
rect 23001 22336 23321 23360
rect 23001 22272 23009 22336
rect 23073 22272 23089 22336
rect 23153 22272 23169 22336
rect 23233 22272 23249 22336
rect 23313 22272 23321 22336
rect 23001 21248 23321 22272
rect 23001 21184 23009 21248
rect 23073 21184 23089 21248
rect 23153 21184 23169 21248
rect 23233 21184 23249 21248
rect 23313 21184 23321 21248
rect 23001 20160 23321 21184
rect 23001 20096 23009 20160
rect 23073 20096 23089 20160
rect 23153 20096 23169 20160
rect 23233 20096 23249 20160
rect 23313 20096 23321 20160
rect 23001 19072 23321 20096
rect 23001 19008 23009 19072
rect 23073 19008 23089 19072
rect 23153 19008 23169 19072
rect 23233 19008 23249 19072
rect 23313 19008 23321 19072
rect 23001 17984 23321 19008
rect 23001 17920 23009 17984
rect 23073 17934 23089 17984
rect 23153 17934 23169 17984
rect 23233 17934 23249 17984
rect 23313 17920 23321 17984
rect 23001 17698 23043 17920
rect 23279 17698 23321 17920
rect 23001 16896 23321 17698
rect 23001 16832 23009 16896
rect 23073 16832 23089 16896
rect 23153 16832 23169 16896
rect 23233 16832 23249 16896
rect 23313 16832 23321 16896
rect 23001 15808 23321 16832
rect 23001 15744 23009 15808
rect 23073 15744 23089 15808
rect 23153 15744 23169 15808
rect 23233 15744 23249 15808
rect 23313 15744 23321 15808
rect 23001 14720 23321 15744
rect 23001 14656 23009 14720
rect 23073 14656 23089 14720
rect 23153 14656 23169 14720
rect 23233 14656 23249 14720
rect 23313 14656 23321 14720
rect 23001 13632 23321 14656
rect 23001 13568 23009 13632
rect 23073 13568 23089 13632
rect 23153 13568 23169 13632
rect 23233 13568 23249 13632
rect 23313 13568 23321 13632
rect 23001 12544 23321 13568
rect 23001 12480 23009 12544
rect 23073 12480 23089 12544
rect 23153 12480 23169 12544
rect 23233 12480 23249 12544
rect 23313 12480 23321 12544
rect 23001 11678 23321 12480
rect 23001 11456 23043 11678
rect 23279 11456 23321 11678
rect 23001 11392 23009 11456
rect 23073 11392 23089 11442
rect 23153 11392 23169 11442
rect 23233 11392 23249 11442
rect 23313 11392 23321 11456
rect 23001 10368 23321 11392
rect 23001 10304 23009 10368
rect 23073 10304 23089 10368
rect 23153 10304 23169 10368
rect 23233 10304 23249 10368
rect 23313 10304 23321 10368
rect 23001 9280 23321 10304
rect 23001 9216 23009 9280
rect 23073 9216 23089 9280
rect 23153 9216 23169 9280
rect 23233 9216 23249 9280
rect 23313 9216 23321 9280
rect 23001 8192 23321 9216
rect 23001 8128 23009 8192
rect 23073 8128 23089 8192
rect 23153 8128 23169 8192
rect 23233 8128 23249 8192
rect 23313 8128 23321 8192
rect 23001 7104 23321 8128
rect 23001 7040 23009 7104
rect 23073 7040 23089 7104
rect 23153 7040 23169 7104
rect 23233 7040 23249 7104
rect 23313 7040 23321 7104
rect 23001 6016 23321 7040
rect 23001 5952 23009 6016
rect 23073 5952 23089 6016
rect 23153 5952 23169 6016
rect 23233 5952 23249 6016
rect 23313 5952 23321 6016
rect 23001 5422 23321 5952
rect 23001 5186 23043 5422
rect 23279 5186 23321 5422
rect 23001 4928 23321 5186
rect 23001 4864 23009 4928
rect 23073 4864 23089 4928
rect 23153 4864 23169 4928
rect 23233 4864 23249 4928
rect 23313 4864 23321 4928
rect 23001 3840 23321 4864
rect 23001 3776 23009 3840
rect 23073 3776 23089 3840
rect 23153 3776 23169 3840
rect 23233 3776 23249 3840
rect 23313 3776 23321 3840
rect 23001 2752 23321 3776
rect 23001 2688 23009 2752
rect 23073 2688 23089 2752
rect 23153 2688 23169 2752
rect 23233 2688 23249 2752
rect 23313 2688 23321 2752
rect 23001 2128 23321 2688
rect 23661 27232 23981 27248
rect 23661 27168 23669 27232
rect 23733 27168 23749 27232
rect 23813 27168 23829 27232
rect 23893 27168 23909 27232
rect 23973 27168 23981 27232
rect 23661 26144 23981 27168
rect 23661 26080 23669 26144
rect 23733 26080 23749 26144
rect 23813 26080 23829 26144
rect 23893 26080 23909 26144
rect 23973 26080 23981 26144
rect 23661 25056 23981 26080
rect 23661 24992 23669 25056
rect 23733 24992 23749 25056
rect 23813 24992 23829 25056
rect 23893 24992 23909 25056
rect 23973 24992 23981 25056
rect 23661 24850 23981 24992
rect 23661 24614 23703 24850
rect 23939 24614 23981 24850
rect 23661 23968 23981 24614
rect 23661 23904 23669 23968
rect 23733 23904 23749 23968
rect 23813 23904 23829 23968
rect 23893 23904 23909 23968
rect 23973 23904 23981 23968
rect 23661 22880 23981 23904
rect 23661 22816 23669 22880
rect 23733 22816 23749 22880
rect 23813 22816 23829 22880
rect 23893 22816 23909 22880
rect 23973 22816 23981 22880
rect 23661 21792 23981 22816
rect 23661 21728 23669 21792
rect 23733 21728 23749 21792
rect 23813 21728 23829 21792
rect 23893 21728 23909 21792
rect 23973 21728 23981 21792
rect 23661 20704 23981 21728
rect 23661 20640 23669 20704
rect 23733 20640 23749 20704
rect 23813 20640 23829 20704
rect 23893 20640 23909 20704
rect 23973 20640 23981 20704
rect 23661 19616 23981 20640
rect 23661 19552 23669 19616
rect 23733 19552 23749 19616
rect 23813 19552 23829 19616
rect 23893 19552 23909 19616
rect 23973 19552 23981 19616
rect 23661 18594 23981 19552
rect 23661 18528 23703 18594
rect 23939 18528 23981 18594
rect 23661 18464 23669 18528
rect 23973 18464 23981 18528
rect 23661 18358 23703 18464
rect 23939 18358 23981 18464
rect 23661 17440 23981 18358
rect 23661 17376 23669 17440
rect 23733 17376 23749 17440
rect 23813 17376 23829 17440
rect 23893 17376 23909 17440
rect 23973 17376 23981 17440
rect 23661 16352 23981 17376
rect 23661 16288 23669 16352
rect 23733 16288 23749 16352
rect 23813 16288 23829 16352
rect 23893 16288 23909 16352
rect 23973 16288 23981 16352
rect 23661 15264 23981 16288
rect 23661 15200 23669 15264
rect 23733 15200 23749 15264
rect 23813 15200 23829 15264
rect 23893 15200 23909 15264
rect 23973 15200 23981 15264
rect 23661 14176 23981 15200
rect 23661 14112 23669 14176
rect 23733 14112 23749 14176
rect 23813 14112 23829 14176
rect 23893 14112 23909 14176
rect 23973 14112 23981 14176
rect 23661 13088 23981 14112
rect 23661 13024 23669 13088
rect 23733 13024 23749 13088
rect 23813 13024 23829 13088
rect 23893 13024 23909 13088
rect 23973 13024 23981 13088
rect 23661 12338 23981 13024
rect 23661 12102 23703 12338
rect 23939 12102 23981 12338
rect 23661 12000 23981 12102
rect 23661 11936 23669 12000
rect 23733 11936 23749 12000
rect 23813 11936 23829 12000
rect 23893 11936 23909 12000
rect 23973 11936 23981 12000
rect 23661 10912 23981 11936
rect 23661 10848 23669 10912
rect 23733 10848 23749 10912
rect 23813 10848 23829 10912
rect 23893 10848 23909 10912
rect 23973 10848 23981 10912
rect 23661 9824 23981 10848
rect 23661 9760 23669 9824
rect 23733 9760 23749 9824
rect 23813 9760 23829 9824
rect 23893 9760 23909 9824
rect 23973 9760 23981 9824
rect 23661 8736 23981 9760
rect 23661 8672 23669 8736
rect 23733 8672 23749 8736
rect 23813 8672 23829 8736
rect 23893 8672 23909 8736
rect 23973 8672 23981 8736
rect 23661 7648 23981 8672
rect 23661 7584 23669 7648
rect 23733 7584 23749 7648
rect 23813 7584 23829 7648
rect 23893 7584 23909 7648
rect 23973 7584 23981 7648
rect 23661 6560 23981 7584
rect 23661 6496 23669 6560
rect 23733 6496 23749 6560
rect 23813 6496 23829 6560
rect 23893 6496 23909 6560
rect 23973 6496 23981 6560
rect 23661 6082 23981 6496
rect 23661 5846 23703 6082
rect 23939 5846 23981 6082
rect 23661 5472 23981 5846
rect 23661 5408 23669 5472
rect 23733 5408 23749 5472
rect 23813 5408 23829 5472
rect 23893 5408 23909 5472
rect 23973 5408 23981 5472
rect 23661 4384 23981 5408
rect 23661 4320 23669 4384
rect 23733 4320 23749 4384
rect 23813 4320 23829 4384
rect 23893 4320 23909 4384
rect 23973 4320 23981 4384
rect 23661 3296 23981 4320
rect 23661 3232 23669 3296
rect 23733 3232 23749 3296
rect 23813 3232 23829 3296
rect 23893 3232 23909 3296
rect 23973 3232 23981 3296
rect 23661 2208 23981 3232
rect 23661 2144 23669 2208
rect 23733 2144 23749 2208
rect 23813 2144 23829 2208
rect 23893 2144 23909 2208
rect 23973 2144 23981 2208
rect 23661 2128 23981 2144
<< via4 >>
rect 4137 23954 4373 24190
rect 4137 17920 4167 17934
rect 4167 17920 4183 17934
rect 4183 17920 4247 17934
rect 4247 17920 4263 17934
rect 4263 17920 4327 17934
rect 4327 17920 4343 17934
rect 4343 17920 4373 17934
rect 4137 17698 4373 17920
rect 4137 11456 4373 11678
rect 4137 11442 4167 11456
rect 4167 11442 4183 11456
rect 4183 11442 4247 11456
rect 4247 11442 4263 11456
rect 4263 11442 4327 11456
rect 4327 11442 4343 11456
rect 4343 11442 4373 11456
rect 4137 5186 4373 5422
rect 4797 24614 5033 24850
rect 10439 23954 10675 24190
rect 4797 18528 5033 18594
rect 4797 18464 4827 18528
rect 4827 18464 4843 18528
rect 4843 18464 4907 18528
rect 4907 18464 4923 18528
rect 4923 18464 4987 18528
rect 4987 18464 5003 18528
rect 5003 18464 5033 18528
rect 4797 18358 5033 18464
rect 10439 17920 10469 17934
rect 10469 17920 10485 17934
rect 10485 17920 10549 17934
rect 10549 17920 10565 17934
rect 10565 17920 10629 17934
rect 10629 17920 10645 17934
rect 10645 17920 10675 17934
rect 10439 17698 10675 17920
rect 4797 12102 5033 12338
rect 10439 11456 10675 11678
rect 10439 11442 10469 11456
rect 10469 11442 10485 11456
rect 10485 11442 10549 11456
rect 10549 11442 10565 11456
rect 10565 11442 10629 11456
rect 10629 11442 10645 11456
rect 10645 11442 10675 11456
rect 4797 5846 5033 6082
rect 10439 5186 10675 5422
rect 11099 24614 11335 24850
rect 11099 18528 11335 18594
rect 11099 18464 11129 18528
rect 11129 18464 11145 18528
rect 11145 18464 11209 18528
rect 11209 18464 11225 18528
rect 11225 18464 11289 18528
rect 11289 18464 11305 18528
rect 11305 18464 11335 18528
rect 11099 18358 11335 18464
rect 11099 12102 11335 12338
rect 11099 5846 11335 6082
rect 16741 23954 16977 24190
rect 16741 17920 16771 17934
rect 16771 17920 16787 17934
rect 16787 17920 16851 17934
rect 16851 17920 16867 17934
rect 16867 17920 16931 17934
rect 16931 17920 16947 17934
rect 16947 17920 16977 17934
rect 16741 17698 16977 17920
rect 16741 11456 16977 11678
rect 16741 11442 16771 11456
rect 16771 11442 16787 11456
rect 16787 11442 16851 11456
rect 16851 11442 16867 11456
rect 16867 11442 16931 11456
rect 16931 11442 16947 11456
rect 16947 11442 16977 11456
rect 16741 5186 16977 5422
rect 17401 24614 17637 24850
rect 17401 18528 17637 18594
rect 17401 18464 17431 18528
rect 17431 18464 17447 18528
rect 17447 18464 17511 18528
rect 17511 18464 17527 18528
rect 17527 18464 17591 18528
rect 17591 18464 17607 18528
rect 17607 18464 17637 18528
rect 17401 18358 17637 18464
rect 17401 12102 17637 12338
rect 17401 5846 17637 6082
rect 23043 23954 23279 24190
rect 23043 17920 23073 17934
rect 23073 17920 23089 17934
rect 23089 17920 23153 17934
rect 23153 17920 23169 17934
rect 23169 17920 23233 17934
rect 23233 17920 23249 17934
rect 23249 17920 23279 17934
rect 23043 17698 23279 17920
rect 23043 11456 23279 11678
rect 23043 11442 23073 11456
rect 23073 11442 23089 11456
rect 23089 11442 23153 11456
rect 23153 11442 23169 11456
rect 23169 11442 23233 11456
rect 23233 11442 23249 11456
rect 23249 11442 23279 11456
rect 23043 5186 23279 5422
rect 23703 24614 23939 24850
rect 23703 18528 23939 18594
rect 23703 18464 23733 18528
rect 23733 18464 23749 18528
rect 23749 18464 23813 18528
rect 23813 18464 23829 18528
rect 23829 18464 23893 18528
rect 23893 18464 23909 18528
rect 23909 18464 23939 18528
rect 23703 18358 23939 18464
rect 23703 12102 23939 12338
rect 23703 5846 23939 6082
<< metal5 >>
rect 1056 24850 26360 24892
rect 1056 24614 4797 24850
rect 5033 24614 11099 24850
rect 11335 24614 17401 24850
rect 17637 24614 23703 24850
rect 23939 24614 26360 24850
rect 1056 24572 26360 24614
rect 1056 24190 26360 24232
rect 1056 23954 4137 24190
rect 4373 23954 10439 24190
rect 10675 23954 16741 24190
rect 16977 23954 23043 24190
rect 23279 23954 26360 24190
rect 1056 23912 26360 23954
rect 1056 18594 26360 18636
rect 1056 18358 4797 18594
rect 5033 18358 11099 18594
rect 11335 18358 17401 18594
rect 17637 18358 23703 18594
rect 23939 18358 26360 18594
rect 1056 18316 26360 18358
rect 1056 17934 26360 17976
rect 1056 17698 4137 17934
rect 4373 17698 10439 17934
rect 10675 17698 16741 17934
rect 16977 17698 23043 17934
rect 23279 17698 26360 17934
rect 1056 17656 26360 17698
rect 1056 12338 26360 12380
rect 1056 12102 4797 12338
rect 5033 12102 11099 12338
rect 11335 12102 17401 12338
rect 17637 12102 23703 12338
rect 23939 12102 26360 12338
rect 1056 12060 26360 12102
rect 1056 11678 26360 11720
rect 1056 11442 4137 11678
rect 4373 11442 10439 11678
rect 10675 11442 16741 11678
rect 16977 11442 23043 11678
rect 23279 11442 26360 11678
rect 1056 11400 26360 11442
rect 1056 6082 26360 6124
rect 1056 5846 4797 6082
rect 5033 5846 11099 6082
rect 11335 5846 17401 6082
rect 17637 5846 23703 6082
rect 23939 5846 26360 6082
rect 1056 5804 26360 5846
rect 1056 5422 26360 5464
rect 1056 5186 4137 5422
rect 4373 5186 10439 5422
rect 10675 5186 16741 5422
rect 16977 5186 23043 5422
rect 23279 5186 26360 5422
rect 1056 5144 26360 5186
use sky130_fd_sc_hd__buf_2  _0676_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _0677_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4600 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0678_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3772 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0679_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3864 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0680_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1683767628
transform 1 0 6164 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0682_
timestamp 1683767628
transform 1 0 6532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0683_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0684_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4508 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0685_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5612 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0686_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 7084 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0687_
timestamp 1683767628
transform 1 0 5704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0688_
timestamp 1683767628
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0689_
timestamp 1683767628
transform 1 0 5152 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0690_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5704 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1683767628
transform 1 0 5888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2760 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0693_
timestamp 1683767628
transform 1 0 3036 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0694_
timestamp 1683767628
transform 1 0 2760 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0695_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0696_
timestamp 1683767628
transform 1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0697_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1656 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0698_
timestamp 1683767628
transform 1 0 3220 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1683767628
transform 1 0 2576 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1683767628
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0701_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4876 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0702_
timestamp 1683767628
transform 1 0 5336 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1683767628
transform 1 0 4968 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1683767628
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0705_
timestamp 1683767628
transform 1 0 4324 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0706_
timestamp 1683767628
transform 1 0 3312 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1683767628
transform 1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0708_
timestamp 1683767628
transform 1 0 3588 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0709_
timestamp 1683767628
transform 1 0 4692 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 1683767628
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0711_
timestamp 1683767628
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0712_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0713_
timestamp 1683767628
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0714_
timestamp 1683767628
transform 1 0 6808 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 1683767628
transform 1 0 7084 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 1683767628
transform 1 0 7360 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0717_
timestamp 1683767628
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0718_
timestamp 1683767628
transform 1 0 6808 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1683767628
transform 1 0 8372 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1683767628
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0721_
timestamp 1683767628
transform 1 0 11684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0722_
timestamp 1683767628
transform 1 0 8924 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0723_
timestamp 1683767628
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0724_
timestamp 1683767628
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0725_
timestamp 1683767628
transform 1 0 7452 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1683767628
transform 1 0 8372 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0727_
timestamp 1683767628
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0728_
timestamp 1683767628
transform 1 0 7084 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1683767628
transform 1 0 8188 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0730_
timestamp 1683767628
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0731_
timestamp 1683767628
transform 1 0 6900 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1683767628
transform 1 0 8004 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0733_
timestamp 1683767628
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0734_
timestamp 1683767628
transform 1 0 5704 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1683767628
transform 1 0 5244 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0736_
timestamp 1683767628
transform 1 0 4968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0737_
timestamp 1683767628
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0738_
timestamp 1683767628
transform 1 0 6348 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 1683767628
transform 1 0 7544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0740_
timestamp 1683767628
transform 1 0 8188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0741_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 11776 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0742_
timestamp 1683767628
transform 1 0 8372 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1683767628
transform 1 0 8464 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0744_
timestamp 1683767628
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0745_
timestamp 1683767628
transform 1 0 5796 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1683767628
transform 1 0 4508 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0747_
timestamp 1683767628
transform 1 0 4048 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0748_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 6348 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0749_
timestamp 1683767628
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0750_
timestamp 1683767628
transform 1 0 6348 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0751_
timestamp 1683767628
transform 1 0 4232 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1683767628
transform 1 0 9752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1683767628
transform 1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1683767628
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0755_
timestamp 1683767628
transform 1 0 5152 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1683767628
transform 1 0 10120 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1683767628
transform 1 0 9384 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0758_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 20700 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1683767628
transform 1 0 22448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0760_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 21160 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0761_
timestamp 1683767628
transform 1 0 23184 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0762_
timestamp 1683767628
transform 1 0 22632 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0763_
timestamp 1683767628
transform 1 0 20700 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0764_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1683767628
transform 1 0 20240 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0766_
timestamp 1683767628
transform 1 0 25024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0767_
timestamp 1683767628
transform 1 0 23644 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0768_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1683767628
transform 1 0 23644 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0770_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 23644 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0771_
timestamp 1683767628
transform 1 0 24380 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1683767628
transform 1 0 24748 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0773_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 24104 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0774_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 20240 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1683767628
transform 1 0 21344 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1683767628
transform 1 0 22724 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0777_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 21804 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0778_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1683767628
transform 1 0 21068 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0780_
timestamp 1683767628
transform 1 0 21804 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0781_
timestamp 1683767628
transform 1 0 22448 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0782_
timestamp 1683767628
transform 1 0 20240 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0783_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0784_
timestamp 1683767628
transform 1 0 21804 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0785_
timestamp 1683767628
transform 1 0 21068 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0786_
timestamp 1683767628
transform 1 0 19504 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1683767628
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0788_
timestamp 1683767628
transform 1 0 20516 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0789_
timestamp 1683767628
transform 1 0 21804 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0790_
timestamp 1683767628
transform 1 0 20700 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0791_
timestamp 1683767628
transform 1 0 20056 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1683767628
transform 1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1683767628
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0794_
timestamp 1683767628
transform 1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1683767628
transform 1 0 21896 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0796_
timestamp 1683767628
transform 1 0 22632 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0797_
timestamp 1683767628
transform 1 0 22632 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0798_
timestamp 1683767628
transform 1 0 21988 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0799_
timestamp 1683767628
transform 1 0 21436 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0800_
timestamp 1683767628
transform 1 0 22080 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0801_
timestamp 1683767628
transform 1 0 22632 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0802_
timestamp 1683767628
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0803_
timestamp 1683767628
transform 1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1683767628
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0805_
timestamp 1683767628
transform 1 0 20332 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0806_
timestamp 1683767628
transform 1 0 20792 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1683767628
transform 1 0 20148 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1683767628
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0809_
timestamp 1683767628
transform 1 0 19320 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0810_
timestamp 1683767628
transform 1 0 19964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0811_
timestamp 1683767628
transform 1 0 20884 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0812_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 20148 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0813_
timestamp 1683767628
transform 1 0 19872 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0814_
timestamp 1683767628
transform 1 0 19228 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0815_
timestamp 1683767628
transform 1 0 15180 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1683767628
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0817_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0818_
timestamp 1683767628
transform 1 0 14076 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0819_
timestamp 1683767628
transform 1 0 14536 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0820_
timestamp 1683767628
transform 1 0 17480 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0821_
timestamp 1683767628
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1683767628
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0823_
timestamp 1683767628
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0824_
timestamp 1683767628
transform 1 0 14536 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0825_
timestamp 1683767628
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0826_
timestamp 1683767628
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0827_
timestamp 1683767628
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0828_
timestamp 1683767628
transform 1 0 13892 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1683767628
transform 1 0 14996 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0830_
timestamp 1683767628
transform 1 0 15180 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0831_
timestamp 1683767628
transform 1 0 14996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1683767628
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1683767628
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0834_
timestamp 1683767628
transform 1 0 15824 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0835_
timestamp 1683767628
transform 1 0 14996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0836_
timestamp 1683767628
transform 1 0 15640 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0837_
timestamp 1683767628
transform 1 0 17388 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0838_
timestamp 1683767628
transform 1 0 16560 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1683767628
transform 1 0 15916 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0840_
timestamp 1683767628
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0841_
timestamp 1683767628
transform 1 0 16652 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0842_
timestamp 1683767628
transform 1 0 15548 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0843_
timestamp 1683767628
transform 1 0 17296 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1683767628
transform 1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0845_
timestamp 1683767628
transform 1 0 17848 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0846_
timestamp 1683767628
transform 1 0 15916 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0847_
timestamp 1683767628
transform 1 0 17020 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0848_
timestamp 1683767628
transform 1 0 17572 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0849_
timestamp 1683767628
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1683767628
transform 1 0 14996 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0851_
timestamp 1683767628
transform 1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1683767628
transform 1 0 15732 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0853_
timestamp 1683767628
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0854_
timestamp 1683767628
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0855_
timestamp 1683767628
transform 1 0 15916 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0856_
timestamp 1683767628
transform 1 0 16560 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0857_
timestamp 1683767628
transform 1 0 16652 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0858_
timestamp 1683767628
transform 1 0 17204 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0859_
timestamp 1683767628
transform 1 0 16376 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0860_
timestamp 1683767628
transform 1 0 17020 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1683767628
transform 1 0 18032 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0862_
timestamp 1683767628
transform 1 0 16652 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0863_
timestamp 1683767628
transform 1 0 17296 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0864_
timestamp 1683767628
transform 1 0 16652 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0865_
timestamp 1683767628
transform 1 0 19964 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1683767628
transform 1 0 18676 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0867_
timestamp 1683767628
transform 1 0 18032 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0868_
timestamp 1683767628
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0869_
timestamp 1683767628
transform 1 0 18584 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0870_
timestamp 1683767628
transform 1 0 18492 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0871_
timestamp 1683767628
transform 1 0 19964 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1683767628
transform 1 0 20792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0873_
timestamp 1683767628
transform 1 0 20976 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0874_
timestamp 1683767628
transform 1 0 19504 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0875_
timestamp 1683767628
transform 1 0 19780 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0876_
timestamp 1683767628
transform 1 0 19872 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0877_
timestamp 1683767628
transform 1 0 19780 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1683767628
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1683767628
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0880_
timestamp 1683767628
transform 1 0 20332 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0881_
timestamp 1683767628
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0882_
timestamp 1683767628
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0883_
timestamp 1683767628
transform 1 0 20240 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0884_
timestamp 1683767628
transform 1 0 19412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1683767628
transform 1 0 20608 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0886_
timestamp 1683767628
transform 1 0 21068 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0887_
timestamp 1683767628
transform 1 0 19412 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0888_
timestamp 1683767628
transform 1 0 21160 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1683767628
transform 1 0 22264 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0890_
timestamp 1683767628
transform 1 0 20608 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0891_
timestamp 1683767628
transform 1 0 20608 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0892_
timestamp 1683767628
transform 1 0 21252 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0893_
timestamp 1683767628
transform 1 0 20976 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0894_
timestamp 1683767628
transform 1 0 21804 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0895_
timestamp 1683767628
transform 1 0 20332 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0896_
timestamp 1683767628
transform 1 0 21068 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0897_
timestamp 1683767628
transform 1 0 20332 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0898_
timestamp 1683767628
transform 1 0 20056 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0899_
timestamp 1683767628
transform 1 0 19688 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1683767628
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0901_
timestamp 1683767628
transform 1 0 21068 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0902_
timestamp 1683767628
transform 1 0 22172 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0903_
timestamp 1683767628
transform 1 0 21528 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0904_
timestamp 1683767628
transform 1 0 21068 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0905_
timestamp 1683767628
transform 1 0 22448 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1683767628
transform 1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1683767628
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1683767628
transform 1 0 22724 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0909_
timestamp 1683767628
transform 1 0 23736 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0910_
timestamp 1683767628
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0911_
timestamp 1683767628
transform 1 0 23184 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0912_
timestamp 1683767628
transform 1 0 22080 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0913_
timestamp 1683767628
transform 1 0 22540 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0914_
timestamp 1683767628
transform 1 0 23092 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0915_
timestamp 1683767628
transform 1 0 19228 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0916_
timestamp 1683767628
transform 1 0 19964 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1683767628
transform 1 0 21160 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0918_
timestamp 1683767628
transform 1 0 20884 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0919_
timestamp 1683767628
transform 1 0 20516 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0920_
timestamp 1683767628
transform 1 0 20240 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0921_
timestamp 1683767628
transform 1 0 20516 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0922_
timestamp 1683767628
transform 1 0 23092 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0923_
timestamp 1683767628
transform 1 0 21252 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0924_
timestamp 1683767628
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0925_
timestamp 1683767628
transform 1 0 21896 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0926_
timestamp 1683767628
transform 1 0 19688 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0927_
timestamp 1683767628
transform 1 0 15272 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1683767628
transform 1 0 16744 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0929_
timestamp 1683767628
transform 1 0 17664 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0930_
timestamp 1683767628
transform 1 0 14628 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0931_
timestamp 1683767628
transform 1 0 15548 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0932_
timestamp 1683767628
transform 1 0 16100 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0933_
timestamp 1683767628
transform 1 0 13248 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1683767628
transform 1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0935_
timestamp 1683767628
transform 1 0 14260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0936_
timestamp 1683767628
transform 1 0 13616 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0937_
timestamp 1683767628
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0938_
timestamp 1683767628
transform 1 0 12880 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0939_
timestamp 1683767628
transform 1 0 13616 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0940_
timestamp 1683767628
transform 1 0 14076 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1683767628
transform 1 0 14720 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0942_
timestamp 1683767628
transform 1 0 14076 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0943_
timestamp 1683767628
transform 1 0 14720 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0944_
timestamp 1683767628
transform 1 0 15364 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1683767628
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0946_
timestamp 1683767628
transform 1 0 15916 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0947_
timestamp 1683767628
transform 1 0 15548 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0948_
timestamp 1683767628
transform 1 0 14904 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0949_
timestamp 1683767628
transform 1 0 17204 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1683767628
transform 1 0 17664 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0951_
timestamp 1683767628
transform 1 0 16468 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0952_
timestamp 1683767628
transform 1 0 16928 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0953_
timestamp 1683767628
transform 1 0 18400 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0954_
timestamp 1683767628
transform 1 0 17020 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0955_
timestamp 1683767628
transform 1 0 9752 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1683767628
transform 1 0 8924 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0957_
timestamp 1683767628
transform 1 0 8372 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1683767628
transform 1 0 9660 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1683767628
transform 1 0 9200 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0960_
timestamp 1683767628
transform 1 0 8372 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0961_
timestamp 1683767628
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1683767628
transform 1 0 11408 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1683767628
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0964_
timestamp 1683767628
transform 1 0 9384 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0965_
timestamp 1683767628
transform 1 0 9660 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0966_
timestamp 1683767628
transform 1 0 9844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0967_
timestamp 1683767628
transform 1 0 9752 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0968_
timestamp 1683767628
transform 1 0 8464 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1683767628
transform 1 0 9200 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0970_
timestamp 1683767628
transform 1 0 9108 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0971_
timestamp 1683767628
transform 1 0 9200 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0972_
timestamp 1683767628
transform 1 0 9752 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1683767628
transform 1 0 8372 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0974_
timestamp 1683767628
transform 1 0 10396 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0975_
timestamp 1683767628
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0976_
timestamp 1683767628
transform 1 0 9476 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0977_
timestamp 1683767628
transform 1 0 7728 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0978_
timestamp 1683767628
transform 1 0 7820 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0979_
timestamp 1683767628
transform 1 0 6532 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0980_
timestamp 1683767628
transform 1 0 7544 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0981_
timestamp 1683767628
transform 1 0 7176 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0982_
timestamp 1683767628
transform 1 0 6808 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _0983_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform -1 0 4876 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0984_
timestamp 1683767628
transform 1 0 5244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0985_
timestamp 1683767628
transform 1 0 14168 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0986_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1683767628
transform 1 0 14536 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0988_
timestamp 1683767628
transform 1 0 13432 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0989_
timestamp 1683767628
transform 1 0 12972 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0990_
timestamp 1683767628
transform 1 0 13616 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0991_
timestamp 1683767628
transform 1 0 12512 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0992_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12880 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 1683767628
transform 1 0 10856 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0994_
timestamp 1683767628
transform 1 0 10580 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0995_
timestamp 1683767628
transform 1 0 14076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1683767628
transform 1 0 21896 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1683767628
transform 1 0 13340 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0998_
timestamp 1683767628
transform 1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0999_
timestamp 1683767628
transform 1 0 14076 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1683767628
transform 1 0 14536 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1001_
timestamp 1683767628
transform 1 0 10580 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1002_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12144 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1003_
timestamp 1683767628
transform 1 0 13892 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1683767628
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1683767628
transform 1 0 14076 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1006_
timestamp 1683767628
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1007_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12236 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1008_
timestamp 1683767628
transform 1 0 13064 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1009_
timestamp 1683767628
transform 1 0 10580 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1010_
timestamp 1683767628
transform 1 0 9844 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1683767628
transform 1 0 9752 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _1012_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10028 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1013_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10396 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1014_
timestamp 1683767628
transform 1 0 12144 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1015_
timestamp 1683767628
transform 1 0 11500 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1683767628
transform 1 0 9936 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1017_
timestamp 1683767628
transform 1 0 13432 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1018_
timestamp 1683767628
transform 1 0 12880 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1019_
timestamp 1683767628
transform 1 0 12144 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1020_
timestamp 1683767628
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1021_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1022_
timestamp 1683767628
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_4  _1023_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10856 0 1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1683767628
transform 1 0 12328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1025_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1683767628
transform 1 0 9016 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1027_
timestamp 1683767628
transform 1 0 8648 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1683767628
transform 1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1683767628
transform 1 0 9752 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1683767628
transform 1 0 10764 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1683767628
transform 1 0 11040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1032_
timestamp 1683767628
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1033_
timestamp 1683767628
transform 1 0 12144 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1683767628
transform 1 0 11960 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1035_
timestamp 1683767628
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1683767628
transform 1 0 11868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1037_
timestamp 1683767628
transform 1 0 11316 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1683767628
transform 1 0 12328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1039_
timestamp 1683767628
transform 1 0 11224 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1040_
timestamp 1683767628
transform 1 0 10028 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1041_
timestamp 1683767628
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1042_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 18308 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1043_
timestamp 1683767628
transform 1 0 13248 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1683767628
transform 1 0 12788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1683767628
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1683767628
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1683767628
transform 1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1683767628
transform 1 0 13064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1683767628
transform 1 0 13708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1683767628
transform 1 0 9752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1683767628
transform 1 0 12788 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1683767628
transform 1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1683767628
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1054_
timestamp 1683767628
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1683767628
transform 1 0 6716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1683767628
transform 1 0 6348 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1683767628
transform 1 0 10304 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1683767628
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1683767628
transform 1 0 6072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1683767628
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1683767628
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1683767628
transform 1 0 10488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1683767628
transform 1 0 10212 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1683767628
transform 1 0 10028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1065_
timestamp 1683767628
transform 1 0 6532 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1683767628
transform 1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1683767628
transform 1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1683767628
transform 1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1683767628
transform 1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1683767628
transform 1 0 2392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1683767628
transform 1 0 2392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1683767628
transform 1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1683767628
transform 1 0 8096 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1683767628
transform 1 0 6900 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1683767628
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1076_
timestamp 1683767628
transform 1 0 4048 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1683767628
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1683767628
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1079_
timestamp 1683767628
transform 1 0 5796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1080_
timestamp 1683767628
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1081_
timestamp 1683767628
transform 1 0 5244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1082_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1683767628
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1084_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5520 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1085_
timestamp 1683767628
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1086_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 4600 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1087_
timestamp 1683767628
transform 1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1088_
timestamp 1683767628
transform 1 0 17480 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1089_
timestamp 1683767628
transform 1 0 18032 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1090_
timestamp 1683767628
transform 1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 1683767628
transform 1 0 13432 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1092_
timestamp 1683767628
transform 1 0 18492 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1093_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 17664 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1094_
timestamp 1683767628
transform 1 0 17848 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1683767628
transform 1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1683767628
transform 1 0 17388 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1097_
timestamp 1683767628
transform 1 0 18584 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1098_
timestamp 1683767628
transform 1 0 9568 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1099_
timestamp 1683767628
transform 1 0 17940 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1100_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 17940 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1101_
timestamp 1683767628
transform 1 0 17296 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1683767628
transform 1 0 17848 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1103_
timestamp 1683767628
transform 1 0 18032 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1104_
timestamp 1683767628
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1683767628
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1106_
timestamp 1683767628
transform 1 0 16744 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1107_
timestamp 1683767628
transform 1 0 12236 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1108_
timestamp 1683767628
transform 1 0 15824 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1109_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 15640 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1110_
timestamp 1683767628
transform 1 0 17848 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1111_
timestamp 1683767628
transform 1 0 16100 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1683767628
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1113_
timestamp 1683767628
transform 1 0 16652 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 1683767628
transform 1 0 10948 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1115_
timestamp 1683767628
transform 1 0 17204 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1683767628
transform 1 0 18308 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1117_
timestamp 1683767628
transform 1 0 17756 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1118_
timestamp 1683767628
transform 1 0 17204 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1119_
timestamp 1683767628
transform 1 0 16836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _1120_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16284 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1121_
timestamp 1683767628
transform 1 0 18860 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1122_
timestamp 1683767628
transform 1 0 17112 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1123_
timestamp 1683767628
transform 1 0 15180 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1124_
timestamp 1683767628
transform 1 0 11500 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1125_
timestamp 1683767628
transform 1 0 16192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1683767628
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1127_
timestamp 1683767628
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1128_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 14352 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _1129_
timestamp 1683767628
transform 1 0 15732 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1130_
timestamp 1683767628
transform 1 0 16192 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1131_
timestamp 1683767628
transform 1 0 15824 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1132_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1133_
timestamp 1683767628
transform 1 0 15732 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1134_
timestamp 1683767628
transform 1 0 17204 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1135_
timestamp 1683767628
transform 1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1136_
timestamp 1683767628
transform 1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1137_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16376 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  _1138_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 15640 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1139_
timestamp 1683767628
transform 1 0 6440 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1140_
timestamp 1683767628
transform 1 0 6624 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1683767628
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1142_
timestamp 1683767628
transform 1 0 23736 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 1683767628
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1683767628
transform 1 0 22540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1683767628
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1683767628
transform 1 0 25300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1683767628
transform 1 0 22448 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1683767628
transform 1 0 22724 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1149_
timestamp 1683767628
transform 1 0 23000 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1683767628
transform 1 0 23736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1683767628
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1683767628
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1153_
timestamp 1683767628
transform 1 0 19412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1683767628
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1155_
timestamp 1683767628
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 1683767628
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1683767628
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1158_
timestamp 1683767628
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1159_
timestamp 1683767628
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1683767628
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1683767628
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1683767628
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1163_
timestamp 1683767628
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1164_
timestamp 1683767628
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1683767628
transform 1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1683767628
transform 1 0 15548 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1167_
timestamp 1683767628
transform 1 0 16192 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1683767628
transform 1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1683767628
transform 1 0 18032 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1683767628
transform 1 0 17756 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1171_
timestamp 1683767628
transform 1 0 19964 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1683767628
transform 1 0 20240 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1683767628
transform 1 0 20700 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1174_
timestamp 1683767628
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1175_
timestamp 1683767628
transform 1 0 23184 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1176_
timestamp 1683767628
transform 1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1177_
timestamp 1683767628
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1683767628
transform 1 0 23920 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1683767628
transform 1 0 23092 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1683767628
transform 1 0 21436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1683767628
transform 1 0 23552 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1683767628
transform 1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1683767628
transform 1 0 23644 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1683767628
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1683767628
transform 1 0 21436 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1186_
timestamp 1683767628
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1683767628
transform 1 0 20424 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1683767628
transform 1 0 20148 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1683767628
transform 1 0 13708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190_
timestamp 1683767628
transform 1 0 14260 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1683767628
transform 1 0 12972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1683767628
transform 1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1683767628
transform 1 0 15272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1194_
timestamp 1683767628
transform 1 0 18952 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1195_
timestamp 1683767628
transform 1 0 19044 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1196_
timestamp 1683767628
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1197_
timestamp 1683767628
transform 1 0 12972 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198_
timestamp 1683767628
transform 1 0 7360 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1199_
timestamp 1683767628
transform 1 0 6808 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1683767628
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1683767628
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1683767628
transform 1 0 6440 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1203_
timestamp 1683767628
transform 1 0 14628 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1204_
timestamp 1683767628
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1683767628
transform 1 0 18860 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1206_
timestamp 1683767628
transform 1 0 17296 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1207_
timestamp 1683767628
transform 1 0 18032 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1208_
timestamp 1683767628
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1209_
timestamp 1683767628
transform 1 0 18216 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1210_
timestamp 1683767628
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1683767628
transform 1 0 13800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1212_
timestamp 1683767628
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1213_
timestamp 1683767628
transform 1 0 18584 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1683767628
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1215_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 16652 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1216_
timestamp 1683767628
transform 1 0 18032 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1217_
timestamp 1683767628
transform 1 0 18676 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1218_
timestamp 1683767628
transform 1 0 19228 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1219_
timestamp 1683767628
transform 1 0 14168 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1683767628
transform 1 0 19228 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1221_
timestamp 1683767628
transform 1 0 14904 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1222_
timestamp 1683767628
transform 1 0 15732 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1223_
timestamp 1683767628
transform 1 0 15732 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1224_
timestamp 1683767628
transform 1 0 15732 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1683767628
transform 1 0 9568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1226_
timestamp 1683767628
transform 1 0 12052 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1227_
timestamp 1683767628
transform 1 0 14996 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1228_
timestamp 1683767628
transform 1 0 17480 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1229_
timestamp 1683767628
transform 1 0 15456 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1230_
timestamp 1683767628
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1231_
timestamp 1683767628
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1232_
timestamp 1683767628
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1233_
timestamp 1683767628
transform 1 0 12972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1234_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1235_
timestamp 1683767628
transform 1 0 13524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1236_
timestamp 1683767628
transform 1 0 12052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1237_
timestamp 1683767628
transform 1 0 17572 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1238_
timestamp 1683767628
transform 1 0 18032 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1239_
timestamp 1683767628
transform 1 0 18676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1240_
timestamp 1683767628
transform 1 0 18584 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1241_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 17848 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1242_
timestamp 1683767628
transform 1 0 11500 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1243_
timestamp 1683767628
transform 1 0 17112 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1244_
timestamp 1683767628
transform 1 0 18124 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1245_
timestamp 1683767628
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1246_
timestamp 1683767628
transform 1 0 18400 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1247_
timestamp 1683767628
transform 1 0 17756 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1248_
timestamp 1683767628
transform 1 0 12880 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1249_
timestamp 1683767628
transform 1 0 12972 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1250_
timestamp 1683767628
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1251_
timestamp 1683767628
transform 1 0 14076 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1252_
timestamp 1683767628
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1253_
timestamp 1683767628
transform 1 0 13524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1254_
timestamp 1683767628
transform 1 0 13156 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1255_
timestamp 1683767628
transform 1 0 13524 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1256_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12696 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1257_
timestamp 1683767628
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1258_
timestamp 1683767628
transform 1 0 13524 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1259_
timestamp 1683767628
transform 1 0 9016 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1683767628
transform 1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1261_
timestamp 1683767628
transform 1 0 11960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1262_
timestamp 1683767628
transform 1 0 7820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1263_
timestamp 1683767628
transform 1 0 8372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1264_
timestamp 1683767628
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1265_
timestamp 1683767628
transform 1 0 9108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1266_
timestamp 1683767628
transform 1 0 10028 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1267_
timestamp 1683767628
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1268_
timestamp 1683767628
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1269_
timestamp 1683767628
transform 1 0 10856 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1270_
timestamp 1683767628
transform 1 0 9660 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1271_
timestamp 1683767628
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1272_
timestamp 1683767628
transform 1 0 10488 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1273_
timestamp 1683767628
transform 1 0 11868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1274_
timestamp 1683767628
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1275_
timestamp 1683767628
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1276_
timestamp 1683767628
transform 1 0 11500 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1277_
timestamp 1683767628
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1278_
timestamp 1683767628
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1279_
timestamp 1683767628
transform 1 0 10396 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1280_
timestamp 1683767628
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1281_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 10764 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1282_
timestamp 1683767628
transform 1 0 10212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1283_
timestamp 1683767628
transform 1 0 12236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1284_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1683767628
transform 1 0 4968 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1286_
timestamp 1683767628
transform 1 0 5796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1683767628
transform 1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1683767628
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1289_
timestamp 1683767628
transform 1 0 6348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1290_
timestamp 1683767628
transform 1 0 7084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1291_
timestamp 1683767628
transform 1 0 7084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1292_
timestamp 1683767628
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1683767628
transform 1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1294_
timestamp 1683767628
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1295_
timestamp 1683767628
transform 1 0 4968 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1296_
timestamp 1683767628
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1297_
timestamp 1683767628
transform 1 0 6992 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1298_
timestamp 1683767628
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1299_
timestamp 1683767628
transform 1 0 7636 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1300_
timestamp 1683767628
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1301_
timestamp 1683767628
transform 1 0 7636 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1683767628
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1303_
timestamp 1683767628
transform 1 0 7636 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1304_
timestamp 1683767628
transform 1 0 8280 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1683767628
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1306_
timestamp 1683767628
transform 1 0 6992 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1307_
timestamp 1683767628
transform 1 0 6440 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1308_
timestamp 1683767628
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1309_
timestamp 1683767628
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1310_
timestamp 1683767628
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1311_
timestamp 1683767628
transform 1 0 4968 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1312_
timestamp 1683767628
transform 1 0 7084 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1313_
timestamp 1683767628
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1314_
timestamp 1683767628
transform 1 0 5428 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1315_
timestamp 1683767628
transform 1 0 5980 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1316_
timestamp 1683767628
transform 1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1317_
timestamp 1683767628
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1318_
timestamp 1683767628
transform 1 0 6624 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1319_
timestamp 1683767628
transform 1 0 4692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1683767628
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1321_
timestamp 1683767628
transform 1 0 5520 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1322_
timestamp 1683767628
transform 1 0 6072 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1323_
timestamp 1683767628
transform 1 0 4416 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1324_
timestamp 1683767628
transform 1 0 5152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1325_
timestamp 1683767628
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1326_
timestamp 1683767628
transform 1 0 4968 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1327_
timestamp 1683767628
transform 1 0 5888 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1328_
timestamp 1683767628
transform 1 0 7360 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1329_
timestamp 1683767628
transform 1 0 6900 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1330_
timestamp 1683767628
transform 1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1331_
timestamp 1683767628
transform 1 0 7084 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1332_
timestamp 1683767628
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1333_
timestamp 1683767628
transform 1 0 3220 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1334_
timestamp 1683767628
transform 1 0 2852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1335_
timestamp 1683767628
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1336_
timestamp 1683767628
transform 1 0 1472 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1337_
timestamp 1683767628
transform 1 0 2116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1338_
timestamp 1683767628
transform 1 0 5980 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1339_
timestamp 1683767628
transform 1 0 4232 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1340_
timestamp 1683767628
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1341_
timestamp 1683767628
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1342_
timestamp 1683767628
transform 1 0 7268 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 1683767628
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1344_
timestamp 1683767628
transform 1 0 6348 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1345_
timestamp 1683767628
transform 1 0 6164 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1346_
timestamp 1683767628
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1347_
timestamp 1683767628
transform 1 0 7084 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1348_
timestamp 1683767628
transform 1 0 7544 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1349_
timestamp 1683767628
transform 1 0 4048 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1350_
timestamp 1683767628
transform 1 0 3772 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1351_
timestamp 1683767628
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1352_
timestamp 1683767628
transform 1 0 4324 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 1683767628
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1354_
timestamp 1683767628
transform 1 0 2668 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1355_
timestamp 1683767628
transform 1 0 3220 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1683767628
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1357_
timestamp 1683767628
transform 1 0 1564 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1358_
timestamp 1683767628
transform 1 0 2300 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1359_
timestamp 1683767628
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1360_
timestamp 1683767628
transform 1 0 2852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1361_
timestamp 1683767628
transform 1 0 2392 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1362_
timestamp 1683767628
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1363_
timestamp 1683767628
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _1364_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 11776 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1365_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 12144 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1366_
timestamp 1683767628
transform 1 0 9200 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1367_
timestamp 1683767628
transform 1 0 12144 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1368_
timestamp 1683767628
transform 1 0 11776 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1369_
timestamp 1683767628
transform 1 0 11868 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1370_
timestamp 1683767628
transform 1 0 9200 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1371_
timestamp 1683767628
transform 1 0 11776 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1372_
timestamp 1683767628
transform 1 0 9660 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1373_
timestamp 1683767628
transform 1 0 9568 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1374_
timestamp 1683767628
transform 1 0 6348 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1375_
timestamp 1683767628
transform 1 0 3772 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1376_
timestamp 1683767628
transform 1 0 9200 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1377_
timestamp 1683767628
transform 1 0 6992 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1378_
timestamp 1683767628
transform 1 0 4416 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1379_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8188 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1380_
timestamp 1683767628
transform 1 0 7544 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1381_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 9292 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1382_
timestamp 1683767628
transform 1 0 9384 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1383_
timestamp 1683767628
transform 1 0 9200 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1384_
timestamp 1683767628
transform 1 0 6992 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1385_
timestamp 1683767628
transform 1 0 1380 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1386_
timestamp 1683767628
transform 1 0 1564 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1387_
timestamp 1683767628
transform 1 0 4140 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1388_
timestamp 1683767628
transform 1 0 1380 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1389_
timestamp 1683767628
transform 1 0 1472 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1390_
timestamp 1683767628
transform 1 0 1380 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1391_
timestamp 1683767628
transform 1 0 5612 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1392_
timestamp 1683767628
transform 1 0 6348 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1393_
timestamp 1683767628
transform 1 0 3588 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1394_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8280 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_2  _1395_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 23092 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1396_
timestamp 1683767628
transform 1 0 20516 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1397_
timestamp 1683767628
transform 1 0 23368 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1398_
timestamp 1683767628
transform 1 0 23552 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1399_
timestamp 1683767628
transform 1 0 20792 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1400_
timestamp 1683767628
transform 1 0 20700 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1401_
timestamp 1683767628
transform 1 0 20792 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1402_
timestamp 1683767628
transform 1 0 22356 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1403_
timestamp 1683767628
transform 1 0 21804 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1404_
timestamp 1683767628
transform 1 0 23000 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1405_
timestamp 1683767628
transform 1 0 21160 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1406_
timestamp 1683767628
transform 1 0 19320 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1407_
timestamp 1683767628
transform 1 0 19228 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1408_
timestamp 1683767628
transform 1 0 18308 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1409_
timestamp 1683767628
transform 1 0 12696 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1410_
timestamp 1683767628
transform 1 0 12880 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1411_
timestamp 1683767628
transform 1 0 12052 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1412_
timestamp 1683767628
transform 1 0 15824 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1413_
timestamp 1683767628
transform 1 0 16468 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1414_
timestamp 1683767628
transform 1 0 16652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1415_
timestamp 1683767628
transform 1 0 14812 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1416_
timestamp 1683767628
transform 1 0 14444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1417_
timestamp 1683767628
transform 1 0 14260 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1418_
timestamp 1683767628
transform 1 0 14076 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1419_
timestamp 1683767628
transform 1 0 16928 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1420_
timestamp 1683767628
transform 1 0 16744 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1421_
timestamp 1683767628
transform 1 0 19228 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1422_
timestamp 1683767628
transform 1 0 18860 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1423_
timestamp 1683767628
transform 1 0 20332 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1424_
timestamp 1683767628
transform 1 0 16652 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1425_
timestamp 1683767628
transform 1 0 21436 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1426_
timestamp 1683767628
transform 1 0 21988 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1427_
timestamp 1683767628
transform 1 0 22080 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1428_
timestamp 1683767628
transform 1 0 21988 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1429_
timestamp 1683767628
transform 1 0 19596 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1430_
timestamp 1683767628
transform 1 0 22172 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1431_
timestamp 1683767628
transform 1 0 22908 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1432_
timestamp 1683767628
transform 1 0 22632 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1433_
timestamp 1683767628
transform 1 0 23000 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1434_
timestamp 1683767628
transform 1 0 19780 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1435_
timestamp 1683767628
transform 1 0 19688 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1436_
timestamp 1683767628
transform 1 0 19412 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1437_
timestamp 1683767628
transform 1 0 12052 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1438_
timestamp 1683767628
transform 1 0 12420 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1439_
timestamp 1683767628
transform 1 0 12052 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1440_
timestamp 1683767628
transform 1 0 11776 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1441_
timestamp 1683767628
transform 1 0 14352 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _1442_
timestamp 1683767628
transform 1 0 17020 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1443_
timestamp 1683767628
transform 1 0 17112 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1444_
timestamp 1683767628
transform 1 0 10212 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1445_
timestamp 1683767628
transform 1 0 12052 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1446_
timestamp 1683767628
transform 1 0 6532 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1447_
timestamp 1683767628
transform 1 0 6348 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1448_
timestamp 1683767628
transform 1 0 10212 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1449_
timestamp 1683767628
transform 1 0 4692 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1450_
timestamp 1683767628
transform 1 0 5612 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1683767628
transform 1 0 11040 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1683767628
transform 1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1683767628
transform 1 0 10396 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1683767628
transform 1 0 11408 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1683767628
transform 1 0 8188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1456_
timestamp 1683767628
transform 1 0 3772 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1683767628
transform 1 0 8096 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1683767628
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1683767628
transform 1 0 5612 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1683767628
transform 1 0 4692 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1461_
timestamp 1683767628
transform 1 0 4324 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1683767628
transform 1 0 9844 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1683767628
transform 1 0 6992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1683767628
transform 1 0 2116 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1683767628
transform 1 0 2116 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1683767628
transform 1 0 3772 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1683767628
transform 1 0 3772 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1683767628
transform 1 0 8096 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1683767628
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1683767628
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1471_
timestamp 1683767628
transform 1 0 2576 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1472_
timestamp 1683767628
transform 1 0 2208 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1473_
timestamp 1683767628
transform 1 0 2208 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1474_
timestamp 1683767628
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform -1 0 3864 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1683767628
transform -1 0 5244 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK_SR pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 6348 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 12604 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CLK_SR
timestamp 1683767628
transform 1 0 5244 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CLK_SR
timestamp 1683767628
transform 1 0 5244 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 5244 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 15640 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 15640 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 10396 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 10396 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 19044 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_Dead_Time_Generator_inst_1.clk
timestamp 1683767628
transform 1 0 18216 0 -1 20672
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_12 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_34
timestamp 1683767628
transform 1 0 4232 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_46 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_52 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 5888 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1683767628
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69
timestamp 1683767628
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1683767628
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1683767628
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1683767628
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_118
timestamp 1683767628
transform 1 0 11960 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_130
timestamp 1683767628
transform 1 0 13064 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_136
timestamp 1683767628
transform 1 0 13616 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1683767628
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 1683767628
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_160
timestamp 1683767628
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1683767628
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1683767628
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1683767628
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1683767628
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_205
timestamp 1683767628
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_212
timestamp 1683767628
transform 1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1683767628
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237
timestamp 1683767628
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_245
timestamp 1683767628
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1683767628
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1683767628
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1683767628
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1683767628
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1683767628
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1683767628
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_63
timestamp 1683767628
transform 1 0 6900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_75
timestamp 1683767628
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_79
timestamp 1683767628
transform 1 0 8372 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_83
timestamp 1683767628
transform 1 0 8740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_95
timestamp 1683767628
transform 1 0 9844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1683767628
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_125
timestamp 1683767628
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_147
timestamp 1683767628
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_159
timestamp 1683767628
transform 1 0 15732 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_190
timestamp 1683767628
transform 1 0 18584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_198
timestamp 1683767628
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_212
timestamp 1683767628
transform 1 0 20608 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_218
timestamp 1683767628
transform 1 0 21160 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_222
timestamp 1683767628
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1683767628
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1683767628
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1683767628
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_261
timestamp 1683767628
transform 1 0 25116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_269
timestamp 1683767628
transform 1 0 25852 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1683767628
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1683767628
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1683767628
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1683767628
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_37
timestamp 1683767628
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_70
timestamp 1683767628
transform 1 0 7544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1683767628
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_117
timestamp 1683767628
transform 1 0 11868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_152
timestamp 1683767628
transform 1 0 15088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_187
timestamp 1683767628
transform 1 0 18308 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_239
timestamp 1683767628
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_246
timestamp 1683767628
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1683767628
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_265
timestamp 1683767628
transform 1 0 25484 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1683767628
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1683767628
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_27
timestamp 1683767628
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1683767628
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_69
timestamp 1683767628
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_92
timestamp 1683767628
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_96
timestamp 1683767628
transform 1 0 9936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_126
timestamp 1683767628
transform 1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_134
timestamp 1683767628
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_138
timestamp 1683767628
transform 1 0 13800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_149
timestamp 1683767628
transform 1 0 14812 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_158
timestamp 1683767628
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_177
timestamp 1683767628
transform 1 0 17388 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_185
timestamp 1683767628
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1683767628
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1683767628
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_241
timestamp 1683767628
transform 1 0 23276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_253
timestamp 1683767628
transform 1 0 24380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_265
timestamp 1683767628
transform 1 0 25484 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1683767628
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1683767628
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1683767628
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1683767628
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_41
timestamp 1683767628
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_45
timestamp 1683767628
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_61
timestamp 1683767628
transform 1 0 6716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_69
timestamp 1683767628
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_74
timestamp 1683767628
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1683767628
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1683767628
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_97
timestamp 1683767628
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_105
timestamp 1683767628
transform 1 0 10764 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_112
timestamp 1683767628
transform 1 0 11408 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1683767628
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_133
timestamp 1683767628
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1683767628
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1683767628
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_156
timestamp 1683767628
transform 1 0 15456 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_173
timestamp 1683767628
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp 1683767628
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1683767628
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1683767628
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1683767628
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1683767628
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_265
timestamp 1683767628
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1683767628
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1683767628
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1683767628
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1683767628
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1683767628
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1683767628
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_75
timestamp 1683767628
transform 1 0 8004 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_87
timestamp 1683767628
transform 1 0 9108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1683767628
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1683767628
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1683767628
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1683767628
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_137
timestamp 1683767628
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_146
timestamp 1683767628
transform 1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_154
timestamp 1683767628
transform 1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_164
timestamp 1683767628
transform 1 0 16192 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_184
timestamp 1683767628
transform 1 0 18032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_196
timestamp 1683767628
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_203
timestamp 1683767628
transform 1 0 19780 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_211
timestamp 1683767628
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1683767628
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1683767628
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_229
timestamp 1683767628
transform 1 0 22172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_233
timestamp 1683767628
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_238
timestamp 1683767628
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_250
timestamp 1683767628
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_262
timestamp 1683767628
transform 1 0 25208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_270
timestamp 1683767628
transform 1 0 25944 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1683767628
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1683767628
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1683767628
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1683767628
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 1683767628
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_76
timestamp 1683767628
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1683767628
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_95
timestamp 1683767628
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_104
timestamp 1683767628
transform 1 0 10672 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_128
timestamp 1683767628
transform 1 0 12880 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_144
timestamp 1683767628
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1683767628
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_186
timestamp 1683767628
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1683767628
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1683767628
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_212
timestamp 1683767628
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_218
timestamp 1683767628
transform 1 0 21160 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_253
timestamp 1683767628
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_257
timestamp 1683767628
transform 1 0 24748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_261
timestamp 1683767628
transform 1 0 25116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_269
timestamp 1683767628
transform 1 0 25852 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1683767628
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1683767628
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1683767628
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_39
timestamp 1683767628
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_71
timestamp 1683767628
transform 1 0 7636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_127
timestamp 1683767628
transform 1 0 12788 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_149
timestamp 1683767628
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1683767628
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_176
timestamp 1683767628
transform 1 0 17296 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1683767628
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_193
timestamp 1683767628
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_220
timestamp 1683767628
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_233
timestamp 1683767628
transform 1 0 22540 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_259
timestamp 1683767628
transform 1 0 24932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1683767628
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1683767628
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1683767628
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_45
timestamp 1683767628
transform 1 0 5244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_66
timestamp 1683767628
transform 1 0 7176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_72
timestamp 1683767628
transform 1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1683767628
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_100
timestamp 1683767628
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_132
timestamp 1683767628
transform 1 0 13248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1683767628
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1683767628
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1683767628
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_165
timestamp 1683767628
transform 1 0 16284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_188
timestamp 1683767628
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_197
timestamp 1683767628
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_222
timestamp 1683767628
transform 1 0 21528 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1683767628
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_245
timestamp 1683767628
transform 1 0 23644 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1683767628
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_265
timestamp 1683767628
transform 1 0 25484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1683767628
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_11
timestamp 1683767628
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_42
timestamp 1683767628
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1683767628
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1683767628
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_69
timestamp 1683767628
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1683767628
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_121
timestamp 1683767628
transform 1 0 12236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_133
timestamp 1683767628
transform 1 0 13340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_145
timestamp 1683767628
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_157
timestamp 1683767628
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1683767628
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1683767628
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_181
timestamp 1683767628
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_197
timestamp 1683767628
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_216
timestamp 1683767628
transform 1 0 20976 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_220
timestamp 1683767628
transform 1 0 21344 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_252
timestamp 1683767628
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_264
timestamp 1683767628
transform 1 0 25392 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_270
timestamp 1683767628
transform 1 0 25944 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1683767628
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_15
timestamp 1683767628
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_40
timestamp 1683767628
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_44
timestamp 1683767628
transform 1 0 5152 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_57
timestamp 1683767628
transform 1 0 6348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_69
timestamp 1683767628
transform 1 0 7452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_73
timestamp 1683767628
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1683767628
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1683767628
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1683767628
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_97
timestamp 1683767628
transform 1 0 10028 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_102
timestamp 1683767628
transform 1 0 10488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_114
timestamp 1683767628
transform 1 0 11592 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_126
timestamp 1683767628
transform 1 0 12696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1683767628
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_149
timestamp 1683767628
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 1683767628
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_203
timestamp 1683767628
transform 1 0 19780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_215
timestamp 1683767628
transform 1 0 20884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_227
timestamp 1683767628
transform 1 0 21988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_241
timestamp 1683767628
transform 1 0 23276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_249
timestamp 1683767628
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1683767628
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_265
timestamp 1683767628
transform 1 0 25484 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_7
timestamp 1683767628
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_19
timestamp 1683767628
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_27
timestamp 1683767628
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_34
timestamp 1683767628
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_38
timestamp 1683767628
transform 1 0 4600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1683767628
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1683767628
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_69
timestamp 1683767628
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_75
timestamp 1683767628
transform 1 0 8004 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_92
timestamp 1683767628
transform 1 0 9568 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_104
timestamp 1683767628
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_125
timestamp 1683767628
transform 1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_142
timestamp 1683767628
transform 1 0 14168 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_154
timestamp 1683767628
transform 1 0 15272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_158
timestamp 1683767628
transform 1 0 15640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1683767628
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_175
timestamp 1683767628
transform 1 0 17204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_181
timestamp 1683767628
transform 1 0 17756 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_191
timestamp 1683767628
transform 1 0 18676 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_203
timestamp 1683767628
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_215
timestamp 1683767628
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1683767628
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_236
timestamp 1683767628
transform 1 0 22816 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_263
timestamp 1683767628
transform 1 0 25300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1683767628
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 1683767628
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_18
timestamp 1683767628
transform 1 0 2760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_35
timestamp 1683767628
transform 1 0 4324 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1683767628
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1683767628
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1683767628
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_85
timestamp 1683767628
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_91
timestamp 1683767628
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_111
timestamp 1683767628
transform 1 0 11316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_126
timestamp 1683767628
transform 1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 1683767628
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_147
timestamp 1683767628
transform 1 0 14628 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_170
timestamp 1683767628
transform 1 0 16744 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_178
timestamp 1683767628
transform 1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1683767628
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_200
timestamp 1683767628
transform 1 0 19504 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_235
timestamp 1683767628
transform 1 0 22724 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_247
timestamp 1683767628
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1683767628
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_256
timestamp 1683767628
transform 1 0 24656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_268
timestamp 1683767628
transform 1 0 25760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1683767628
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_28
timestamp 1683767628
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1683767628
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_76
timestamp 1683767628
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_103
timestamp 1683767628
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1683767628
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_125
timestamp 1683767628
transform 1 0 12604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_147
timestamp 1683767628
transform 1 0 14628 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_157
timestamp 1683767628
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1683767628
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_201
timestamp 1683767628
transform 1 0 19596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1683767628
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_232
timestamp 1683767628
transform 1 0 22448 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_267
timestamp 1683767628
transform 1 0 25668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_3
timestamp 1683767628
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1683767628
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_41
timestamp 1683767628
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1683767628
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1683767628
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1683767628
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_89
timestamp 1683767628
transform 1 0 9292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_101
timestamp 1683767628
transform 1 0 10396 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_109
timestamp 1683767628
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_119
timestamp 1683767628
transform 1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_129
timestamp 1683767628
transform 1 0 12972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1683767628
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_147
timestamp 1683767628
transform 1 0 14628 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_155
timestamp 1683767628
transform 1 0 15364 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_168
timestamp 1683767628
transform 1 0 16560 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_173
timestamp 1683767628
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_183
timestamp 1683767628
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_187
timestamp 1683767628
transform 1 0 18308 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 1683767628
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_202
timestamp 1683767628
transform 1 0 19688 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_239
timestamp 1683767628
transform 1 0 23092 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_266
timestamp 1683767628
transform 1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_270
timestamp 1683767628
transform 1 0 25944 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1683767628
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_11
timestamp 1683767628
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_19
timestamp 1683767628
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_31
timestamp 1683767628
transform 1 0 3956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_43
timestamp 1683767628
transform 1 0 5060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_47
timestamp 1683767628
transform 1 0 5428 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_62
timestamp 1683767628
transform 1 0 6808 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_74
timestamp 1683767628
transform 1 0 7912 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_88
timestamp 1683767628
transform 1 0 9200 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_100
timestamp 1683767628
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_117
timestamp 1683767628
transform 1 0 11868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_129
timestamp 1683767628
transform 1 0 12972 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_141
timestamp 1683767628
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_153
timestamp 1683767628
transform 1 0 15180 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_162
timestamp 1683767628
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1683767628
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_181
timestamp 1683767628
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_185
timestamp 1683767628
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_202
timestamp 1683767628
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_214
timestamp 1683767628
transform 1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_231
timestamp 1683767628
transform 1 0 22356 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_243
timestamp 1683767628
transform 1 0 23460 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_262
timestamp 1683767628
transform 1 0 25208 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_270
timestamp 1683767628
transform 1 0 25944 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1683767628
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1683767628
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1683767628
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_32
timestamp 1683767628
transform 1 0 4048 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_64
timestamp 1683767628
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_85
timestamp 1683767628
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_109
timestamp 1683767628
transform 1 0 11132 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_122
timestamp 1683767628
transform 1 0 12328 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_134
timestamp 1683767628
transform 1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1683767628
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_152
timestamp 1683767628
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_161
timestamp 1683767628
transform 1 0 15916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_173
timestamp 1683767628
transform 1 0 17020 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1683767628
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1683767628
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_204
timestamp 1683767628
transform 1 0 19872 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_212
timestamp 1683767628
transform 1 0 20608 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_238
timestamp 1683767628
transform 1 0 23000 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_244
timestamp 1683767628
transform 1 0 23552 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_257
timestamp 1683767628
transform 1 0 24748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_269
timestamp 1683767628
transform 1 0 25852 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1683767628
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_22
timestamp 1683767628
transform 1 0 3128 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_28
timestamp 1683767628
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_32
timestamp 1683767628
transform 1 0 4048 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_41
timestamp 1683767628
transform 1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1683767628
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_64
timestamp 1683767628
transform 1 0 6992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_79
timestamp 1683767628
transform 1 0 8372 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_119
timestamp 1683767628
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_133
timestamp 1683767628
transform 1 0 13340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_141
timestamp 1683767628
transform 1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1683767628
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1683767628
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_195
timestamp 1683767628
transform 1 0 19044 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_207
timestamp 1683767628
transform 1 0 20148 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1683767628
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_237
timestamp 1683767628
transform 1 0 22908 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_268
timestamp 1683767628
transform 1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_3
timestamp 1683767628
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1683767628
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 1683767628
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_50
timestamp 1683767628
transform 1 0 5704 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1683767628
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_97
timestamp 1683767628
transform 1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1683767628
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1683767628
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1683767628
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_154
timestamp 1683767628
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_172
timestamp 1683767628
transform 1 0 16928 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_176
timestamp 1683767628
transform 1 0 17296 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_188
timestamp 1683767628
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1683767628
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_209
timestamp 1683767628
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_236
timestamp 1683767628
transform 1 0 22816 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 1683767628
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_256
timestamp 1683767628
transform 1 0 24656 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_268
timestamp 1683767628
transform 1 0 25760 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_9
timestamp 1683767628
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_27
timestamp 1683767628
transform 1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1683767628
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_84
timestamp 1683767628
transform 1 0 8832 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_90
timestamp 1683767628
transform 1 0 9384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1683767628
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1683767628
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_149
timestamp 1683767628
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_153
timestamp 1683767628
transform 1 0 15180 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_157
timestamp 1683767628
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1683767628
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_183
timestamp 1683767628
transform 1 0 17940 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_189
timestamp 1683767628
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_197
timestamp 1683767628
transform 1 0 19228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_209
timestamp 1683767628
transform 1 0 20332 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_225
timestamp 1683767628
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_241
timestamp 1683767628
transform 1 0 23276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_253
timestamp 1683767628
transform 1 0 24380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_265
timestamp 1683767628
transform 1 0 25484 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1683767628
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1683767628
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1683767628
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_66
timestamp 1683767628
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_73
timestamp 1683767628
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1683767628
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1683767628
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_97
timestamp 1683767628
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_108
timestamp 1683767628
transform 1 0 11040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_118
timestamp 1683767628
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_125
timestamp 1683767628
transform 1 0 12604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_130
timestamp 1683767628
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1683767628
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_212
timestamp 1683767628
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_234
timestamp 1683767628
transform 1 0 22632 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_246
timestamp 1683767628
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1683767628
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_265
timestamp 1683767628
transform 1 0 25484 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1683767628
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1683767628
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_27
timestamp 1683767628
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_33
timestamp 1683767628
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_40
timestamp 1683767628
transform 1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_46
timestamp 1683767628
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1683767628
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_62
timestamp 1683767628
transform 1 0 6808 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_71
timestamp 1683767628
transform 1 0 7636 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_79
timestamp 1683767628
transform 1 0 8372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_99
timestamp 1683767628
transform 1 0 10212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1683767628
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1683767628
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_140
timestamp 1683767628
transform 1 0 13984 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_152
timestamp 1683767628
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1683767628
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1683767628
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_178
timestamp 1683767628
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_191
timestamp 1683767628
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_214
timestamp 1683767628
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1683767628
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1683767628
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1683767628
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1683767628
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_261
timestamp 1683767628
transform 1 0 25116 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_269
timestamp 1683767628
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1683767628
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1683767628
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1683767628
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_29
timestamp 1683767628
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_44
timestamp 1683767628
transform 1 0 5152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_48
timestamp 1683767628
transform 1 0 5520 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_52
timestamp 1683767628
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_56
timestamp 1683767628
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_60
timestamp 1683767628
transform 1 0 6624 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_116
timestamp 1683767628
transform 1 0 11776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_149
timestamp 1683767628
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_156
timestamp 1683767628
transform 1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1683767628
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_220
timestamp 1683767628
transform 1 0 21344 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_232
timestamp 1683767628
transform 1 0 22448 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_244
timestamp 1683767628
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1683767628
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_265
timestamp 1683767628
transform 1 0 25484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_23
timestamp 1683767628
transform 1 0 3220 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_31
timestamp 1683767628
transform 1 0 3956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_77
timestamp 1683767628
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1683767628
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_121
timestamp 1683767628
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_165
timestamp 1683767628
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_174
timestamp 1683767628
transform 1 0 17112 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_180
timestamp 1683767628
transform 1 0 17664 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_187
timestamp 1683767628
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_196
timestamp 1683767628
transform 1 0 19136 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_204
timestamp 1683767628
transform 1 0 19872 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_211
timestamp 1683767628
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_216
timestamp 1683767628
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1683767628
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1683767628
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1683767628
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_261
timestamp 1683767628
transform 1 0 25116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_269
timestamp 1683767628
transform 1 0 25852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1683767628
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_25
timestamp 1683767628
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_38
timestamp 1683767628
transform 1 0 4600 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_44
timestamp 1683767628
transform 1 0 5152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1683767628
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1683767628
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_96
timestamp 1683767628
transform 1 0 9936 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_103
timestamp 1683767628
transform 1 0 10580 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_115
timestamp 1683767628
transform 1 0 11684 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_120
timestamp 1683767628
transform 1 0 12144 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_132
timestamp 1683767628
transform 1 0 13248 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1683767628
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1683767628
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_153
timestamp 1683767628
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_160
timestamp 1683767628
transform 1 0 15824 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_182
timestamp 1683767628
transform 1 0 17848 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_187
timestamp 1683767628
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1683767628
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_203
timestamp 1683767628
transform 1 0 19780 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_230
timestamp 1683767628
transform 1 0 22264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_242
timestamp 1683767628
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1683767628
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1683767628
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_265
timestamp 1683767628
transform 1 0 25484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1683767628
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_23
timestamp 1683767628
transform 1 0 3220 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_33
timestamp 1683767628
transform 1 0 4140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_41
timestamp 1683767628
transform 1 0 4876 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1683767628
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1683767628
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_66
timestamp 1683767628
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_80
timestamp 1683767628
transform 1 0 8464 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_92
timestamp 1683767628
transform 1 0 9568 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_98
timestamp 1683767628
transform 1 0 10120 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_103
timestamp 1683767628
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1683767628
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 1683767628
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_119
timestamp 1683767628
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_127
timestamp 1683767628
transform 1 0 12788 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_135
timestamp 1683767628
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_147
timestamp 1683767628
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_159
timestamp 1683767628
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1683767628
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1683767628
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1683767628
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_229
timestamp 1683767628
transform 1 0 22172 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_241
timestamp 1683767628
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_253
timestamp 1683767628
transform 1 0 24380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_265
timestamp 1683767628
transform 1 0 25484 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_6
timestamp 1683767628
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_18
timestamp 1683767628
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1683767628
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_29
timestamp 1683767628
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_57
timestamp 1683767628
transform 1 0 6348 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_63
timestamp 1683767628
transform 1 0 6900 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_88
timestamp 1683767628
transform 1 0 9200 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_144
timestamp 1683767628
transform 1 0 14352 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_156
timestamp 1683767628
transform 1 0 15456 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_168
timestamp 1683767628
transform 1 0 16560 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_174
timestamp 1683767628
transform 1 0 17112 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_178
timestamp 1683767628
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_190
timestamp 1683767628
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_197
timestamp 1683767628
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_214
timestamp 1683767628
transform 1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_220
timestamp 1683767628
transform 1 0 21344 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1683767628
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1683767628
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1683767628
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_265
timestamp 1683767628
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1683767628
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_17
timestamp 1683767628
transform 1 0 2668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_29
timestamp 1683767628
transform 1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_35
timestamp 1683767628
transform 1 0 4324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_69
timestamp 1683767628
transform 1 0 7452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_91
timestamp 1683767628
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 1683767628
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_120
timestamp 1683767628
transform 1 0 12144 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_132
timestamp 1683767628
transform 1 0 13248 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_138
timestamp 1683767628
transform 1 0 13800 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_144
timestamp 1683767628
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_152
timestamp 1683767628
transform 1 0 15088 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_164
timestamp 1683767628
transform 1 0 16192 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_190
timestamp 1683767628
transform 1 0 18584 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_198
timestamp 1683767628
transform 1 0 19320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_206
timestamp 1683767628
transform 1 0 20056 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1683767628
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_225
timestamp 1683767628
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_250
timestamp 1683767628
transform 1 0 24104 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_262
timestamp 1683767628
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_266
timestamp 1683767628
transform 1 0 25576 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1683767628
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_69
timestamp 1683767628
transform 1 0 7452 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_88
timestamp 1683767628
transform 1 0 9200 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_127
timestamp 1683767628
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1683767628
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_149
timestamp 1683767628
transform 1 0 14812 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_161
timestamp 1683767628
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_169
timestamp 1683767628
transform 1 0 16652 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_177
timestamp 1683767628
transform 1 0 17388 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_186
timestamp 1683767628
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1683767628
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_197
timestamp 1683767628
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_205
timestamp 1683767628
transform 1 0 19964 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_211
timestamp 1683767628
transform 1 0 20516 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_224
timestamp 1683767628
transform 1 0 21712 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_232
timestamp 1683767628
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_237
timestamp 1683767628
transform 1 0 22908 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_246
timestamp 1683767628
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1683767628
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_265
timestamp 1683767628
transform 1 0 25484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1683767628
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_14
timestamp 1683767628
transform 1 0 2392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_25
timestamp 1683767628
transform 1 0 3404 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_89
timestamp 1683767628
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_101
timestamp 1683767628
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_125
timestamp 1683767628
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_150
timestamp 1683767628
transform 1 0 14904 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_162
timestamp 1683767628
transform 1 0 16008 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_186
timestamp 1683767628
transform 1 0 18216 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_198
timestamp 1683767628
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_202
timestamp 1683767628
transform 1 0 19688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_208
timestamp 1683767628
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1683767628
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1683767628
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1683767628
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_249
timestamp 1683767628
transform 1 0 24012 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_257
timestamp 1683767628
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_263
timestamp 1683767628
transform 1 0 25300 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 1683767628
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_11
timestamp 1683767628
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_16
timestamp 1683767628
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1683767628
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_41
timestamp 1683767628
transform 1 0 4876 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_72
timestamp 1683767628
transform 1 0 7728 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1683767628
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_93
timestamp 1683767628
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_103
timestamp 1683767628
transform 1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1683767628
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_121
timestamp 1683767628
transform 1 0 12236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1683767628
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_149
timestamp 1683767628
transform 1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_157
timestamp 1683767628
transform 1 0 15548 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_192
timestamp 1683767628
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1683767628
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_226
timestamp 1683767628
transform 1 0 21896 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1683767628
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1683767628
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_265
timestamp 1683767628
transform 1 0 25484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_28
timestamp 1683767628
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_41
timestamp 1683767628
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1683767628
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_60
timestamp 1683767628
transform 1 0 6624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_72
timestamp 1683767628
transform 1 0 7728 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_78
timestamp 1683767628
transform 1 0 8280 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_82
timestamp 1683767628
transform 1 0 8648 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_88
timestamp 1683767628
transform 1 0 9200 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_141
timestamp 1683767628
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_153
timestamp 1683767628
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_157
timestamp 1683767628
transform 1 0 15548 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_198
timestamp 1683767628
transform 1 0 19320 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1683767628
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_233
timestamp 1683767628
transform 1 0 22540 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_242
timestamp 1683767628
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_254
timestamp 1683767628
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_266
timestamp 1683767628
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_270
timestamp 1683767628
transform 1 0 25944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_3
timestamp 1683767628
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_11
timestamp 1683767628
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_17
timestamp 1683767628
transform 1 0 2668 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_40
timestamp 1683767628
transform 1 0 4784 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_48
timestamp 1683767628
transform 1 0 5520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_70
timestamp 1683767628
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_74
timestamp 1683767628
transform 1 0 7912 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1683767628
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_113
timestamp 1683767628
transform 1 0 11500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_121
timestamp 1683767628
transform 1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_130
timestamp 1683767628
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1683767628
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_144
timestamp 1683767628
transform 1 0 14352 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_156
timestamp 1683767628
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_172
timestamp 1683767628
transform 1 0 16928 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_180
timestamp 1683767628
transform 1 0 17664 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_187
timestamp 1683767628
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1683767628
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_203
timestamp 1683767628
transform 1 0 19780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_213
timestamp 1683767628
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_225
timestamp 1683767628
transform 1 0 21804 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1683767628
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1683767628
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_265
timestamp 1683767628
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1683767628
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_15
timestamp 1683767628
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_26
timestamp 1683767628
transform 1 0 3496 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_32
timestamp 1683767628
transform 1 0 4048 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_49
timestamp 1683767628
transform 1 0 5612 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1683767628
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1683767628
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_70
timestamp 1683767628
transform 1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_76
timestamp 1683767628
transform 1 0 8096 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 1683767628
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1683767628
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1683767628
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_125
timestamp 1683767628
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_132
timestamp 1683767628
transform 1 0 13248 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_139
timestamp 1683767628
transform 1 0 13892 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_151
timestamp 1683767628
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1683767628
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_175
timestamp 1683767628
transform 1 0 17204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_181
timestamp 1683767628
transform 1 0 17756 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_206
timestamp 1683767628
transform 1 0 20056 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1683767628
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1683767628
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_258
timestamp 1683767628
transform 1 0 24840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_270
timestamp 1683767628
transform 1 0 25944 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_13
timestamp 1683767628
transform 1 0 2300 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_79
timestamp 1683767628
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1683767628
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_94
timestamp 1683767628
transform 1 0 9752 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_100
timestamp 1683767628
transform 1 0 10304 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_121
timestamp 1683767628
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_132
timestamp 1683767628
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_141
timestamp 1683767628
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_146
timestamp 1683767628
transform 1 0 14536 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_158
timestamp 1683767628
transform 1 0 15640 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_169
timestamp 1683767628
transform 1 0 16652 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_177
timestamp 1683767628
transform 1 0 17388 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_183
timestamp 1683767628
transform 1 0 17940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1683767628
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_197
timestamp 1683767628
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_224
timestamp 1683767628
transform 1 0 21712 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_236
timestamp 1683767628
transform 1 0 22816 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_240
timestamp 1683767628
transform 1 0 23184 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_244
timestamp 1683767628
transform 1 0 23552 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_250
timestamp 1683767628
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_261
timestamp 1683767628
transform 1 0 25116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_269
timestamp 1683767628
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 1683767628
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_77
timestamp 1683767628
transform 1 0 8188 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_88
timestamp 1683767628
transform 1 0 9200 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1683767628
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_121
timestamp 1683767628
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1683767628
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_169
timestamp 1683767628
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_173
timestamp 1683767628
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_181
timestamp 1683767628
transform 1 0 17756 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_191
timestamp 1683767628
transform 1 0 18676 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_203
timestamp 1683767628
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_215
timestamp 1683767628
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1683767628
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1683767628
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1683767628
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1683767628
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_261
timestamp 1683767628
transform 1 0 25116 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_267
timestamp 1683767628
transform 1 0 25668 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1683767628
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1683767628
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1683767628
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_33
timestamp 1683767628
transform 1 0 4140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_45
timestamp 1683767628
transform 1 0 5244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_49
timestamp 1683767628
transform 1 0 5612 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_56
timestamp 1683767628
transform 1 0 6256 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_62
timestamp 1683767628
transform 1 0 6808 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_66
timestamp 1683767628
transform 1 0 7176 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_78
timestamp 1683767628
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_88
timestamp 1683767628
transform 1 0 9200 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_111
timestamp 1683767628
transform 1 0 11316 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_156
timestamp 1683767628
transform 1 0 15456 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_170
timestamp 1683767628
transform 1 0 16744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_174
timestamp 1683767628
transform 1 0 17112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1683767628
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 1683767628
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_201
timestamp 1683767628
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1683767628
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_224
timestamp 1683767628
transform 1 0 21712 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_236
timestamp 1683767628
transform 1 0 22816 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_244
timestamp 1683767628
transform 1 0 23552 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_248
timestamp 1683767628
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1683767628
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_265
timestamp 1683767628
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1683767628
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1683767628
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_27
timestamp 1683767628
transform 1 0 3588 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_31
timestamp 1683767628
transform 1 0 3956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_35
timestamp 1683767628
transform 1 0 4324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_46
timestamp 1683767628
transform 1 0 5336 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1683767628
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1683767628
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_81
timestamp 1683767628
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_89
timestamp 1683767628
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_97
timestamp 1683767628
transform 1 0 10028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_105
timestamp 1683767628
transform 1 0 10764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_118
timestamp 1683767628
transform 1 0 11960 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_139
timestamp 1683767628
transform 1 0 13892 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_151
timestamp 1683767628
transform 1 0 14996 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1683767628
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_176
timestamp 1683767628
transform 1 0 17296 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_196
timestamp 1683767628
transform 1 0 19136 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_225
timestamp 1683767628
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_255
timestamp 1683767628
transform 1 0 24564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_267
timestamp 1683767628
transform 1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1683767628
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1683767628
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1683767628
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_60
timestamp 1683767628
transform 1 0 6624 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_72
timestamp 1683767628
transform 1 0 7728 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_85
timestamp 1683767628
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_93
timestamp 1683767628
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1683767628
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1683767628
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1683767628
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1683767628
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1683767628
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1683767628
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1683767628
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_165
timestamp 1683767628
transform 1 0 16284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_169
timestamp 1683767628
transform 1 0 16652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_177
timestamp 1683767628
transform 1 0 17388 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1683767628
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1683767628
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_197
timestamp 1683767628
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_227
timestamp 1683767628
transform 1 0 21988 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1683767628
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1683767628
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_265
timestamp 1683767628
transform 1 0 25484 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1683767628
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1683767628
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_27
timestamp 1683767628
transform 1 0 3588 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_30
timestamp 1683767628
transform 1 0 3864 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_41
timestamp 1683767628
transform 1 0 4876 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_49
timestamp 1683767628
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1683767628
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_57
timestamp 1683767628
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_61
timestamp 1683767628
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_69
timestamp 1683767628
transform 1 0 7452 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_87
timestamp 1683767628
transform 1 0 9108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_108
timestamp 1683767628
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_116
timestamp 1683767628
transform 1 0 11776 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_128
timestamp 1683767628
transform 1 0 12880 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_132
timestamp 1683767628
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_146
timestamp 1683767628
transform 1 0 14536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_152
timestamp 1683767628
transform 1 0 15088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_156
timestamp 1683767628
transform 1 0 15456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 1683767628
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1683767628
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1683767628
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1683767628
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_205
timestamp 1683767628
transform 1 0 19964 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1683767628
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_225
timestamp 1683767628
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_259
timestamp 1683767628
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1683767628
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1683767628
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1683767628
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1683767628
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_41
timestamp 1683767628
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_78
timestamp 1683767628
transform 1 0 8280 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_98
timestamp 1683767628
transform 1 0 10120 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_168
timestamp 1683767628
transform 1 0 16560 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_174
timestamp 1683767628
transform 1 0 17112 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_182
timestamp 1683767628
transform 1 0 17848 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 1683767628
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1683767628
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_209
timestamp 1683767628
transform 1 0 20332 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_221
timestamp 1683767628
transform 1 0 21436 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_229
timestamp 1683767628
transform 1 0 22172 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_235
timestamp 1683767628
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1683767628
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_256
timestamp 1683767628
transform 1 0 24656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_268
timestamp 1683767628
transform 1 0 25760 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1683767628
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1683767628
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1683767628
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1683767628
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_54
timestamp 1683767628
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_57
timestamp 1683767628
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_78
timestamp 1683767628
transform 1 0 8280 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_82
timestamp 1683767628
transform 1 0 8648 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_98
timestamp 1683767628
transform 1 0 10120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1683767628
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1683767628
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_125
timestamp 1683767628
transform 1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_132
timestamp 1683767628
transform 1 0 13248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_153
timestamp 1683767628
transform 1 0 15180 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_158
timestamp 1683767628
transform 1 0 15640 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_162
timestamp 1683767628
transform 1 0 16008 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_198
timestamp 1683767628
transform 1 0 19320 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_225
timestamp 1683767628
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_236
timestamp 1683767628
transform 1 0 22816 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_248
timestamp 1683767628
transform 1 0 23920 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_260
timestamp 1683767628
transform 1 0 25024 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_268
timestamp 1683767628
transform 1 0 25760 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1683767628
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1683767628
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1683767628
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_29
timestamp 1683767628
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_37
timestamp 1683767628
transform 1 0 4508 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_65
timestamp 1683767628
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_71
timestamp 1683767628
transform 1 0 7636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1683767628
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_85
timestamp 1683767628
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_122
timestamp 1683767628
transform 1 0 12328 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_128
timestamp 1683767628
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1683767628
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1683767628
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_145
timestamp 1683767628
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_149
timestamp 1683767628
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_163
timestamp 1683767628
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1683767628
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_197
timestamp 1683767628
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_226
timestamp 1683767628
transform 1 0 21896 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_230
timestamp 1683767628
transform 1 0 22264 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_247
timestamp 1683767628
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1683767628
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_261
timestamp 1683767628
transform 1 0 25116 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_267
timestamp 1683767628
transform 1 0 25668 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1683767628
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1683767628
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1683767628
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1683767628
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1683767628
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1683767628
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_104
timestamp 1683767628
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_140
timestamp 1683767628
transform 1 0 13984 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_169
timestamp 1683767628
transform 1 0 16652 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_197
timestamp 1683767628
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_201
timestamp 1683767628
transform 1 0 19596 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1683767628
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_225
timestamp 1683767628
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_250
timestamp 1683767628
transform 1 0 24104 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_262
timestamp 1683767628
transform 1 0 25208 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_270
timestamp 1683767628
transform 1 0 25944 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1683767628
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1683767628
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1683767628
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1683767628
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1683767628
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_53
timestamp 1683767628
transform 1 0 5980 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_80
timestamp 1683767628
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_85
timestamp 1683767628
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1683767628
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_109
timestamp 1683767628
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_117
timestamp 1683767628
transform 1 0 11868 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1683767628
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_153
timestamp 1683767628
transform 1 0 15180 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_157
timestamp 1683767628
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_166
timestamp 1683767628
transform 1 0 16376 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_172
timestamp 1683767628
transform 1 0 16928 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_185
timestamp 1683767628
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1683767628
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 1683767628
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_205
timestamp 1683767628
transform 1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_213
timestamp 1683767628
transform 1 0 20700 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_225
timestamp 1683767628
transform 1 0 21804 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_237
timestamp 1683767628
transform 1 0 22908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_249
timestamp 1683767628
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1683767628
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_265
timestamp 1683767628
transform 1 0 25484 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_6
timestamp 1683767628
transform 1 0 1656 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_18
timestamp 1683767628
transform 1 0 2760 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_26
timestamp 1683767628
transform 1 0 3496 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_35
timestamp 1683767628
transform 1 0 4324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_47
timestamp 1683767628
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1683767628
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_57
timestamp 1683767628
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_65
timestamp 1683767628
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_72
timestamp 1683767628
transform 1 0 7728 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_85
timestamp 1683767628
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_97
timestamp 1683767628
transform 1 0 10028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_109
timestamp 1683767628
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_113
timestamp 1683767628
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_121
timestamp 1683767628
transform 1 0 12236 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_133
timestamp 1683767628
transform 1 0 13340 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_139
timestamp 1683767628
transform 1 0 13892 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_141
timestamp 1683767628
transform 1 0 14076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_153
timestamp 1683767628
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_160
timestamp 1683767628
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1683767628
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1683767628
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_193
timestamp 1683767628
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_197
timestamp 1683767628
transform 1 0 19228 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1683767628
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1683767628
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1683767628
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1683767628
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_237
timestamp 1683767628
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_247
timestamp 1683767628
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_251
timestamp 1683767628
transform 1 0 24196 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_253
timestamp 1683767628
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_265
timestamp 1683767628
transform 1 0 25484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold6
timestamp 1683767628
transform 1 0 9292 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1683767628
transform 1 0 9292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold8
timestamp 1683767628
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1683767628
transform 1 0 10304 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1683767628
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1683767628
transform 1 0 11316 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold12
timestamp 1683767628
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1683767628
transform 1 0 7360 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold14
timestamp 1683767628
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1683767628
transform 1 0 10120 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1683767628
transform 1 0 12512 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1683767628
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1683767628
transform 1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1683767628
transform 1 0 8096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1683767628
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1683767628
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1683767628
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1683767628
transform 1 0 15640 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1683767628
transform 1 0 12696 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1683767628
transform 1 0 9568 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1683767628
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1683767628
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1683767628
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1683767628
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1683767628
transform 1 0 12512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1683767628
transform 1 0 4968 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1683767628
transform 1 0 14444 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1683767628
transform 1 0 17480 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1683767628
transform 1 0 14260 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1683767628
transform 1 0 22540 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1683767628
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold37
timestamp 1683767628
transform 1 0 14536 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  hold38
timestamp 1683767628
transform 1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1683767628
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold41
timestamp 1683767628
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1683767628
transform 1 0 2668 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1683767628
transform 1 0 16560 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1683767628
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1683767628
transform 1 0 11960 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1683767628
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1683767628
transform 1 0 5244 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1683767628
transform 1 0 21988 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1683767628
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1683767628
transform 1 0 25024 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1683767628
transform 1 0 5612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1683767628
transform 1 0 17572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1683767628
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1683767628
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1683767628
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1683767628
transform 1 0 22356 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1683767628
transform 1 0 14904 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1683767628
transform 1 0 15640 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1683767628
transform 1 0 11040 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1683767628
transform 1 0 11224 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1683767628
transform 1 0 4140 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1683767628
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1683767628
transform 1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1683767628
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1683767628
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1683767628
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1683767628
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1683767628
transform 1 0 25760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1683767628
transform 1 0 25760 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1683767628
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1683767628
transform 1 0 15548 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1683767628
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1683767628
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1683767628
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1683767628
transform 1 0 25760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1683767628
transform 1 0 7176 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1683767628
transform 1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1683767628
transform 1 0 25484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1683767628
transform 1 0 23276 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1683767628
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1683767628
transform 1 0 25668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1683767628
transform 1 0 19412 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1683767628
transform 1 0 25484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1683767628
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1683767628
transform 1 0 3772 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output25 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 1380 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1683767628
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1683767628
transform -1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1683767628
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1683767628
transform -1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1683767628
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1683767628
transform -1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1683767628
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1683767628
transform -1 0 26312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1683767628
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1683767628
transform -1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1683767628
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1683767628
transform -1 0 26312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1683767628
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1683767628
transform -1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1683767628
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1683767628
transform -1 0 26312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1683767628
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1683767628
transform -1 0 26312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1683767628
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1683767628
transform -1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1683767628
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1683767628
transform -1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1683767628
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1683767628
transform -1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1683767628
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1683767628
transform -1 0 26312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1683767628
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1683767628
transform -1 0 26312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1683767628
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1683767628
transform -1 0 26312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1683767628
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1683767628
transform -1 0 26312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1683767628
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1683767628
transform -1 0 26312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1683767628
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1683767628
transform -1 0 26312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1683767628
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1683767628
transform -1 0 26312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1683767628
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1683767628
transform -1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1683767628
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1683767628
transform -1 0 26312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1683767628
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1683767628
transform -1 0 26312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1683767628
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1683767628
transform -1 0 26312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1683767628
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1683767628
transform -1 0 26312 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1683767628
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1683767628
transform -1 0 26312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1683767628
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1683767628
transform -1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1683767628
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1683767628
transform -1 0 26312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1683767628
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1683767628
transform -1 0 26312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1683767628
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1683767628
transform -1 0 26312 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1683767628
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1683767628
transform -1 0 26312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1683767628
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1683767628
transform -1 0 26312 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1683767628
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1683767628
transform -1 0 26312 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1683767628
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1683767628
transform -1 0 26312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1683767628
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1683767628
transform -1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1683767628
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1683767628
transform -1 0 26312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1683767628
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1683767628
transform -1 0 26312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1683767628
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1683767628
transform -1 0 26312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1683767628
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1683767628
transform -1 0 26312 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1683767628
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1683767628
transform -1 0 26312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1683767628
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1683767628
transform -1 0 26312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1683767628
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1683767628
transform -1 0 26312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1683767628
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1683767628
transform -1 0 26312 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1683767628
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1683767628
transform -1 0 26312 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1683767628
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1683767628
transform -1 0 26312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1683767628
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1683767628
transform -1 0 26312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1683767628
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1683767628
transform -1 0 26312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1683767628
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1683767628
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1683767628
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1683767628
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1683767628
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1683767628
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1683767628
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1683767628
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1683767628
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1683767628
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1683767628
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1683767628
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1683767628
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1683767628
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1683767628
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1683767628
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1683767628
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1683767628
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1683767628
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1683767628
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1683767628
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1683767628
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1683767628
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1683767628
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1683767628
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1683767628
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1683767628
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1683767628
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1683767628
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1683767628
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1683767628
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1683767628
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1683767628
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1683767628
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1683767628
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1683767628
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1683767628
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1683767628
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1683767628
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1683767628
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1683767628
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1683767628
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1683767628
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1683767628
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1683767628
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1683767628
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1683767628
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1683767628
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1683767628
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1683767628
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1683767628
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1683767628
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1683767628
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1683767628
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1683767628
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1683767628
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1683767628
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1683767628
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1683767628
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1683767628
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1683767628
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1683767628
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1683767628
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1683767628
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1683767628
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1683767628
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1683767628
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1683767628
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1683767628
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1683767628
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1683767628
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1683767628
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1683767628
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1683767628
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1683767628
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1683767628
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1683767628
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1683767628
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1683767628
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1683767628
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1683767628
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1683767628
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1683767628
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1683767628
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1683767628
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1683767628
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1683767628
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1683767628
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1683767628
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1683767628
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1683767628
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1683767628
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1683767628
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1683767628
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1683767628
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1683767628
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1683767628
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1683767628
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1683767628
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1683767628
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1683767628
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1683767628
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1683767628
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1683767628
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1683767628
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1683767628
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1683767628
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1683767628
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1683767628
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1683767628
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1683767628
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1683767628
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1683767628
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1683767628
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1683767628
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1683767628
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1683767628
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1683767628
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1683767628
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1683767628
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1683767628
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1683767628
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1683767628
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1683767628
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1683767628
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1683767628
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1683767628
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1683767628
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1683767628
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1683767628
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1683767628
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1683767628
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1683767628
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1683767628
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1683767628
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1683767628
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1683767628
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1683767628
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1683767628
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1683767628
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1683767628
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1683767628
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1683767628
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1683767628
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1683767628
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1683767628
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1683767628
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1683767628
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1683767628
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1683767628
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1683767628
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1683767628
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1683767628
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1683767628
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1683767628
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1683767628
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1683767628
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1683767628
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1683767628
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1683767628
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1683767628
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1683767628
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1683767628
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1683767628
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1683767628
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1683767628
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1683767628
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1683767628
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1683767628
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1683767628
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1683767628
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1683767628
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1683767628
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1683767628
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1683767628
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1683767628
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1683767628
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1683767628
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1683767628
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1683767628
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1683767628
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1683767628
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1683767628
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1683767628
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1683767628
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1683767628
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1683767628
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1683767628
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1683767628
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1683767628
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1683767628
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1683767628
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1683767628
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1683767628
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1683767628
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1683767628
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1683767628
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1683767628
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1683767628
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1683767628
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1683767628
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1683767628
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1683767628
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1683767628
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1683767628
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1683767628
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1683767628
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1683767628
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1683767628
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1683767628
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1683767628
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1683767628
transform 1 0 13984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1683767628
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1683767628
transform 1 0 19136 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1683767628
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1683767628
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 CLK_EXT
port 0 nsew signal input
flabel metal2 s 27066 28825 27122 29625 0 FreeSans 224 90 0 0 CLK_PLL
port 1 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 CLK_SR
port 2 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 Data_SR
port 3 nsew signal input
flabel metal2 s 7102 28825 7158 29625 0 FreeSans 224 90 0 0 NMOS1_PS1
port 4 nsew signal tristate
flabel metal2 s 11610 28825 11666 29625 0 FreeSans 224 90 0 0 NMOS1_PS2
port 5 nsew signal tristate
flabel metal3 s 26681 8168 27481 8288 0 FreeSans 480 0 0 0 NMOS2_PS1
port 6 nsew signal tristate
flabel metal2 s 23202 28825 23258 29625 0 FreeSans 224 90 0 0 NMOS2_PS2
port 7 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 NMOS_PS3
port 8 nsew signal tristate
flabel metal3 s 26681 17008 27481 17128 0 FreeSans 480 0 0 0 PMOS1_PS1
port 9 nsew signal tristate
flabel metal2 s 19338 28825 19394 29625 0 FreeSans 224 90 0 0 PMOS1_PS2
port 10 nsew signal tristate
flabel metal3 s 26681 8 27481 128 0 FreeSans 480 0 0 0 PMOS2_PS1
port 11 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 PMOS2_PS2
port 12 nsew signal tristate
flabel metal2 s 3238 28825 3294 29625 0 FreeSans 224 90 0 0 PMOS_PS3
port 13 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 RST
port 14 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 SIGNAL_OUTPUT
port 15 nsew signal tristate
flabel metal4 s 4755 2128 5075 27248 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 11057 2128 11377 27248 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 17359 2128 17679 27248 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 23661 2128 23981 27248 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 5804 26360 6124 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 12060 26360 12380 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 18316 26360 18636 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 24572 26360 24892 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 4095 2128 4415 27248 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 10397 2128 10717 27248 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 16699 2128 17019 27248 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 23001 2128 23321 27248 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 5144 26360 5464 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 11400 26360 11720 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 17656 26360 17976 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 23912 26360 24232 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 d1[0]
port 18 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 d1[1]
port 19 nsew signal input
flabel metal3 s 26681 4088 27481 4208 0 FreeSans 480 0 0 0 d1[2]
port 20 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 d1[3]
port 21 nsew signal input
flabel metal3 s 26681 21088 27481 21208 0 FreeSans 480 0 0 0 d1[4]
port 22 nsew signal input
flabel metal3 s 26681 25168 27481 25288 0 FreeSans 480 0 0 0 d1[5]
port 23 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 d2[0]
port 24 nsew signal input
flabel metal2 s 15474 28825 15530 29625 0 FreeSans 224 90 0 0 d2[1]
port 25 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 d2[2]
port 26 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 d2[3]
port 27 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 d2[4]
port 28 nsew signal input
flabel metal3 s 26681 12928 27481 13048 0 FreeSans 480 0 0 0 d2[5]
port 29 nsew signal input
rlabel metal1 13708 27200 13708 27200 0 VGND
rlabel metal1 13708 26656 13708 26656 0 VPWR
rlabel metal3 2200 4148 2200 4148 0 CLK_EXT
rlabel via2 5198 23749 5198 23749 0 CLK_PLL
rlabel metal1 4830 18326 4830 18326 0 CLK_SR
rlabel metal3 1050 8228 1050 8228 0 Data_SR
rlabel via2 12650 15045 12650 15045 0 Dead_Time_Generator_inst_1.clk
rlabel metal1 10442 7888 10442 7888 0 Dead_Time_Generator_inst_1.count_dt\[0\]
rlabel metal2 8326 6018 8326 6018 0 Dead_Time_Generator_inst_1.count_dt\[1\]
rlabel metal2 12006 4828 12006 4828 0 Dead_Time_Generator_inst_1.count_dt\[2\]
rlabel metal1 10948 6222 10948 6222 0 Dead_Time_Generator_inst_1.count_dt\[3\]
rlabel metal2 9614 7004 9614 7004 0 Dead_Time_Generator_inst_1.count_dt\[4\]
rlabel metal1 5612 17510 5612 17510 0 Dead_Time_Generator_inst_1.dt\[0\]
rlabel metal2 5658 8041 5658 8041 0 Dead_Time_Generator_inst_1.dt\[1\]
rlabel metal1 9706 5713 9706 5713 0 Dead_Time_Generator_inst_1.dt\[2\]
rlabel metal1 6532 12750 6532 12750 0 Dead_Time_Generator_inst_1.dt\[3\]
rlabel metal1 4416 14382 4416 14382 0 Dead_Time_Generator_inst_1.dt\[4\]
rlabel metal1 11500 10030 11500 10030 0 Dead_Time_Generator_inst_1.go
rlabel metal1 7774 5168 7774 5168 0 Dead_Time_Generator_inst_2.count_dt\[0\]
rlabel metal1 7866 3434 7866 3434 0 Dead_Time_Generator_inst_2.count_dt\[1\]
rlabel metal2 7130 6256 7130 6256 0 Dead_Time_Generator_inst_2.count_dt\[2\]
rlabel metal2 5842 3808 5842 3808 0 Dead_Time_Generator_inst_2.count_dt\[3\]
rlabel metal1 5014 6392 5014 6392 0 Dead_Time_Generator_inst_2.count_dt\[4\]
rlabel metal2 9522 9078 9522 9078 0 Dead_Time_Generator_inst_2.go
rlabel metal2 7682 11373 7682 11373 0 Dead_Time_Generator_inst_3.count_dt\[0\]
rlabel metal1 6256 13294 6256 13294 0 Dead_Time_Generator_inst_3.count_dt\[1\]
rlabel metal2 3542 13056 3542 13056 0 Dead_Time_Generator_inst_3.count_dt\[2\]
rlabel metal1 5612 13430 5612 13430 0 Dead_Time_Generator_inst_3.count_dt\[3\]
rlabel metal2 5198 13124 5198 13124 0 Dead_Time_Generator_inst_3.count_dt\[4\]
rlabel metal1 8694 11322 8694 11322 0 Dead_Time_Generator_inst_3.go
rlabel metal1 6348 10710 6348 10710 0 Dead_Time_Generator_inst_4.count_dt\[0\]
rlabel metal1 5566 7854 5566 7854 0 Dead_Time_Generator_inst_4.count_dt\[1\]
rlabel metal1 4692 8534 4692 8534 0 Dead_Time_Generator_inst_4.count_dt\[2\]
rlabel metal2 3450 9146 3450 9146 0 Dead_Time_Generator_inst_4.count_dt\[3\]
rlabel metal1 3818 8840 3818 8840 0 Dead_Time_Generator_inst_4.count_dt\[4\]
rlabel metal1 11454 9554 11454 9554 0 Dead_Time_Generator_inst_4.go
rlabel metal1 7268 27098 7268 27098 0 NMOS1_PS1
rlabel metal2 13938 16048 13938 16048 0 NMOS1_PS1_prev
rlabel metal1 11868 27098 11868 27098 0 NMOS1_PS2
rlabel metal1 13716 19482 13716 19482 0 NMOS1_PS2_prev
rlabel metal2 25898 8279 25898 8279 0 NMOS2_PS1
rlabel metal1 13984 16762 13984 16762 0 NMOS2_PS1_prev
rlabel metal2 23506 27319 23506 27319 0 NMOS2_PS2
rlabel metal2 12926 15810 12926 15810 0 NMOS2_PS2_prev
rlabel metal2 20010 1520 20010 1520 0 NMOS_PS3
rlabel via2 25898 17051 25898 17051 0 PMOS1_PS1
rlabel metal1 13961 12954 13961 12954 0 PMOS1_PS1_prev
rlabel metal1 19504 27098 19504 27098 0 PMOS1_PS2
rlabel via1 13593 12410 13593 12410 0 PMOS1_PS2_prev
rlabel metal1 25254 2278 25254 2278 0 PMOS2_PS1
rlabel metal1 10925 11866 10925 11866 0 PMOS2_PS1_prev
rlabel metal3 1142 12308 1142 12308 0 PMOS2_PS2
rlabel via1 11063 11322 11063 11322 0 PMOS2_PS2_prev
rlabel metal1 3634 27098 3634 27098 0 PMOS_PS3
rlabel metal2 23874 1027 23874 1027 0 RST
rlabel metal2 46 1554 46 1554 0 SIGNAL_OUTPUT
rlabel metal2 9982 20128 9982 20128 0 Shift_Register_Inst.data_out\[10\]
rlabel metal1 10718 16014 10718 16014 0 Shift_Register_Inst.data_out\[11\]
rlabel metal1 8740 16762 8740 16762 0 Shift_Register_Inst.data_out\[12\]
rlabel metal1 11500 13362 11500 13362 0 Shift_Register_Inst.data_out\[13\]
rlabel metal1 5612 23290 5612 23290 0 Shift_Register_Inst.data_out\[14\]
rlabel metal1 7866 15130 7866 15130 0 Shift_Register_Inst.data_out\[15\]
rlabel metal1 13248 18054 13248 18054 0 Shift_Register_Inst.data_out\[16\]
rlabel metal1 12788 18258 12788 18258 0 Shift_Register_Inst.data_out\[17\]
rlabel metal1 14812 10030 14812 10030 0 Shift_Register_Inst.data_out\[5\]
rlabel metal2 15318 9962 15318 9962 0 Shift_Register_Inst.data_out\[6\]
rlabel metal1 17066 22032 17066 22032 0 Shift_Register_Inst.data_out\[7\]
rlabel metal1 15042 21658 15042 21658 0 Shift_Register_Inst.data_out\[8\]
rlabel metal2 9338 17816 9338 17816 0 Shift_Register_Inst.data_out\[9\]
rlabel metal1 2852 20434 2852 20434 0 Shift_Register_Inst.shift_state\[0\]
rlabel metal2 2990 19652 2990 19652 0 Shift_Register_Inst.shift_state\[1\]
rlabel metal2 7314 20434 7314 20434 0 Shift_Register_Inst.shift_state\[2\]
rlabel metal1 7590 20910 7590 20910 0 Shift_Register_Inst.shift_state\[3\]
rlabel metal1 5474 21454 5474 21454 0 Shift_Register_Inst.shift_state\[4\]
rlabel metal1 21068 9554 21068 9554 0 Signal_Generator_1_0phase_inst.count\[0\]
rlabel metal2 21022 9248 21022 9248 0 Signal_Generator_1_0phase_inst.count\[1\]
rlabel metal1 19182 9996 19182 9996 0 Signal_Generator_1_0phase_inst.count\[2\]
rlabel metal1 20838 9452 20838 9452 0 Signal_Generator_1_0phase_inst.count\[3\]
rlabel metal1 20378 11322 20378 11322 0 Signal_Generator_1_0phase_inst.count\[4\]
rlabel metal1 22494 13158 22494 13158 0 Signal_Generator_1_0phase_inst.count\[5\]
rlabel metal1 21298 12818 21298 12818 0 Signal_Generator_1_0phase_inst.direction
rlabel metal1 14260 5134 14260 5134 0 Signal_Generator_1_180phase_inst.count\[0\]
rlabel metal1 15295 6970 15295 6970 0 Signal_Generator_1_180phase_inst.count\[1\]
rlabel metal1 16054 6358 16054 6358 0 Signal_Generator_1_180phase_inst.count\[2\]
rlabel metal1 18377 6970 18377 6970 0 Signal_Generator_1_180phase_inst.count\[3\]
rlabel metal1 18170 5882 18170 5882 0 Signal_Generator_1_180phase_inst.count\[4\]
rlabel metal1 16905 9146 16905 9146 0 Signal_Generator_1_180phase_inst.count\[5\]
rlabel metal1 17480 6154 17480 6154 0 Signal_Generator_1_180phase_inst.direction
rlabel metal1 16606 13260 16606 13260 0 Signal_Generator_1_270phase_inst.count\[0\]
rlabel metal1 16974 12716 16974 12716 0 Signal_Generator_1_270phase_inst.count\[1\]
rlabel metal1 17304 9622 17304 9622 0 Signal_Generator_1_270phase_inst.count\[2\]
rlabel viali 17810 9622 17810 9622 0 Signal_Generator_1_270phase_inst.count\[3\]
rlabel metal1 20102 13294 20102 13294 0 Signal_Generator_1_270phase_inst.count\[4\]
rlabel metal2 20378 13600 20378 13600 0 Signal_Generator_1_270phase_inst.count\[5\]
rlabel metal1 17940 14382 17940 14382 0 Signal_Generator_1_270phase_inst.direction
rlabel metal1 18400 6766 18400 6766 0 Signal_Generator_1_90phase_inst.count\[0\]
rlabel metal1 22356 6290 22356 6290 0 Signal_Generator_1_90phase_inst.count\[1\]
rlabel metal1 19090 6970 19090 6970 0 Signal_Generator_1_90phase_inst.count\[2\]
rlabel metal2 19090 6494 19090 6494 0 Signal_Generator_1_90phase_inst.count\[3\]
rlabel metal1 19596 4998 19596 4998 0 Signal_Generator_1_90phase_inst.count\[4\]
rlabel metal1 20378 4556 20378 4556 0 Signal_Generator_1_90phase_inst.count\[5\]
rlabel metal1 21206 4522 21206 4522 0 Signal_Generator_1_90phase_inst.direction
rlabel metal1 17526 17578 17526 17578 0 Signal_Generator_2_0phase_inst.count\[0\]
rlabel metal1 19228 19346 19228 19346 0 Signal_Generator_2_0phase_inst.count\[1\]
rlabel metal1 20470 17204 20470 17204 0 Signal_Generator_2_0phase_inst.count\[2\]
rlabel metal1 18699 18666 18699 18666 0 Signal_Generator_2_0phase_inst.count\[3\]
rlabel metal1 17894 20468 17894 20468 0 Signal_Generator_2_0phase_inst.count\[4\]
rlabel metal2 21390 21284 21390 21284 0 Signal_Generator_2_0phase_inst.count\[5\]
rlabel metal2 21022 15844 21022 15844 0 Signal_Generator_2_0phase_inst.direction
rlabel metal1 14398 21998 14398 21998 0 Signal_Generator_2_180phase_inst.count\[0\]
rlabel metal1 15594 24242 15594 24242 0 Signal_Generator_2_180phase_inst.count\[1\]
rlabel metal1 16422 23494 16422 23494 0 Signal_Generator_2_180phase_inst.count\[2\]
rlabel metal2 16376 24242 16376 24242 0 Signal_Generator_2_180phase_inst.count\[3\]
rlabel metal1 18124 24786 18124 24786 0 Signal_Generator_2_180phase_inst.count\[4\]
rlabel metal1 16974 24378 16974 24378 0 Signal_Generator_2_180phase_inst.count\[5\]
rlabel metal1 16790 25942 16790 25942 0 Signal_Generator_2_180phase_inst.direction
rlabel metal1 13846 21998 13846 21998 0 Signal_Generator_2_270phase_inst.count\[0\]
rlabel metal1 9338 25296 9338 25296 0 Signal_Generator_2_270phase_inst.count\[1\]
rlabel via2 10810 23188 10810 23188 0 Signal_Generator_2_270phase_inst.count\[2\]
rlabel metal1 12052 24038 12052 24038 0 Signal_Generator_2_270phase_inst.count\[3\]
rlabel metal2 13018 22950 13018 22950 0 Signal_Generator_2_270phase_inst.count\[4\]
rlabel metal1 8694 23664 8694 23664 0 Signal_Generator_2_270phase_inst.count\[5\]
rlabel metal1 9706 26248 9706 26248 0 Signal_Generator_2_270phase_inst.direction
rlabel metal2 14122 21250 14122 21250 0 Signal_Generator_2_90phase_inst.count\[0\]
rlabel metal1 18078 21352 18078 21352 0 Signal_Generator_2_90phase_inst.count\[1\]
rlabel metal1 18630 21998 18630 21998 0 Signal_Generator_2_90phase_inst.count\[2\]
rlabel metal1 19780 21998 19780 21998 0 Signal_Generator_2_90phase_inst.count\[3\]
rlabel metal1 19734 24174 19734 24174 0 Signal_Generator_2_90phase_inst.count\[4\]
rlabel metal1 20378 21862 20378 21862 0 Signal_Generator_2_90phase_inst.count\[5\]
rlabel metal1 20470 24854 20470 24854 0 Signal_Generator_2_90phase_inst.direction
rlabel metal2 12466 14620 12466 14620 0 _0000_
rlabel metal1 12098 15130 12098 15130 0 _0001_
rlabel metal2 12466 16082 12466 16082 0 _0002_
rlabel metal1 12052 13974 12052 13974 0 _0003_
rlabel metal1 10994 12274 10994 12274 0 _0004_
rlabel metal2 11638 11764 11638 11764 0 _0005_
rlabel metal1 9246 10778 9246 10778 0 _0006_
rlabel metal1 10028 12682 10028 12682 0 _0007_
rlabel metal1 20608 8874 20608 8874 0 _0008_
rlabel metal1 23644 11254 23644 11254 0 _0009_
rlabel metal1 24012 9622 24012 9622 0 _0010_
rlabel metal2 21114 10268 21114 10268 0 _0011_
rlabel metal2 20930 12002 20930 12002 0 _0012_
rlabel metal2 21114 13090 21114 13090 0 _0013_
rlabel metal2 24058 11492 24058 11492 0 _0014_
rlabel metal2 13294 6460 13294 6460 0 _0015_
rlabel metal2 12466 3604 12466 3604 0 _0016_
rlabel metal1 16008 3502 16008 3502 0 _0017_
rlabel metal1 16744 6766 16744 6766 0 _0018_
rlabel metal2 17066 3434 17066 3434 0 _0019_
rlabel metal1 15410 5338 15410 5338 0 _0020_
rlabel via1 14030 3366 14030 3366 0 _0021_
rlabel metal2 14582 11934 14582 11934 0 _0022_
rlabel metal1 14398 13192 14398 13192 0 _0023_
rlabel metal2 17802 15844 17802 15844 0 _0024_
rlabel metal1 17204 13158 17204 13158 0 _0025_
rlabel metal1 19550 14280 19550 14280 0 _0026_
rlabel metal1 18906 13362 18906 13362 0 _0027_
rlabel metal1 15824 14246 15824 14246 0 _0028_
rlabel metal1 21896 7310 21896 7310 0 _0029_
rlabel metal1 23230 6290 23230 6290 0 _0030_
rlabel metal2 22678 3740 22678 3740 0 _0031_
rlabel metal1 20240 6426 20240 6426 0 _0032_
rlabel metal2 19642 3740 19642 3740 0 _0033_
rlabel metal1 18952 4046 18952 4046 0 _0034_
rlabel metal2 22770 5508 22770 5508 0 _0035_
rlabel metal1 16698 17238 16698 17238 0 _0036_
rlabel metal2 21850 16218 21850 16218 0 _0037_
rlabel metal2 22310 17374 22310 17374 0 _0038_
rlabel metal1 22241 18666 22241 18666 0 _0039_
rlabel metal1 22310 19720 22310 19720 0 _0040_
rlabel metal1 20010 20026 20010 20026 0 _0041_
rlabel metal1 20792 15470 20792 15470 0 _0042_
rlabel metal1 13432 21454 13432 21454 0 _0043_
rlabel metal2 12466 24412 12466 24412 0 _0044_
rlabel metal1 14076 24650 14076 24650 0 _0045_
rlabel metal2 15502 25636 15502 25636 0 _0046_
rlabel metal1 17066 24922 17066 24922 0 _0047_
rlabel metal1 17388 25262 17388 25262 0 _0048_
rlabel metal1 12880 25398 12880 25398 0 _0049_
rlabel metal1 11960 21930 11960 21930 0 _0050_
rlabel metal1 8372 26418 8372 26418 0 _0051_
rlabel metal1 6670 25976 6670 25976 0 _0052_
rlabel metal1 10534 24072 10534 24072 0 _0053_
rlabel metal1 7038 24378 7038 24378 0 _0054_
rlabel metal1 6854 23800 6854 23800 0 _0055_
rlabel metal1 10396 25330 10396 25330 0 _0056_
rlabel metal1 23368 20434 23368 20434 0 _0057_
rlabel metal1 23000 22610 23000 22610 0 _0058_
rlabel metal1 23460 23698 23460 23698 0 _0059_
rlabel metal1 20286 22542 20286 22542 0 _0060_
rlabel metal1 20240 24922 20240 24922 0 _0061_
rlabel metal2 19734 25058 19734 25058 0 _0062_
rlabel metal1 22540 24378 22540 24378 0 _0063_
rlabel metal2 12926 13022 12926 13022 0 _0064_
rlabel metal1 13945 16490 13945 16490 0 _0065_
rlabel metal1 10626 11723 10626 11723 0 _0066_
rlabel metal1 13570 14423 13570 14423 0 _0067_
rlabel metal2 13202 12002 13202 12002 0 _0068_
rlabel metal1 13623 13974 13623 13974 0 _0069_
rlabel metal2 9936 11628 9936 11628 0 _0070_
rlabel metal2 12834 19550 12834 19550 0 _0071_
rlabel metal1 11224 18938 11224 18938 0 _0072_
rlabel metal1 11369 19414 11369 19414 0 _0073_
rlabel metal1 6992 14586 6992 14586 0 _0074_
rlabel metal1 5895 23018 5895 23018 0 _0075_
rlabel metal2 10258 14824 10258 14824 0 _0076_
rlabel metal1 8793 16490 8793 16490 0 _0077_
rlabel metal2 6210 16898 6210 16898 0 _0078_
rlabel metal2 9246 20264 9246 20264 0 _0079_
rlabel metal1 9016 17510 9016 17510 0 _0080_
rlabel metal1 10863 21590 10863 21590 0 _0081_
rlabel metal2 10350 22168 10350 22168 0 _0082_
rlabel metal2 10166 15198 10166 15198 0 _0083_
rlabel metal1 8188 15334 8188 15334 0 _0084_
rlabel metal2 2806 15470 2806 15470 0 _0085_
rlabel metal2 2990 15674 2990 15674 0 _0086_
rlabel metal2 5750 14824 5750 14824 0 _0087_
rlabel metal1 2484 17306 2484 17306 0 _0088_
rlabel metal2 2530 21352 2530 21352 0 _0089_
rlabel metal2 2806 19142 2806 19142 0 _0090_
rlabel metal1 7505 20842 7505 20842 0 _0091_
rlabel metal2 7130 21726 7130 21726 0 _0092_
rlabel metal2 3542 21352 3542 21352 0 _0093_
rlabel metal2 24518 11934 24518 11934 0 _0094_
rlabel metal2 22678 8738 22678 8738 0 _0095_
rlabel metal2 24426 8670 24426 8670 0 _0096_
rlabel metal2 25438 9758 25438 9758 0 _0097_
rlabel metal1 22494 9146 22494 9146 0 _0098_
rlabel metal1 22586 12614 22586 12614 0 _0099_
rlabel metal2 23138 13090 23138 13090 0 _0100_
rlabel metal2 23598 6120 23598 6120 0 _0101_
rlabel metal1 22494 6834 22494 6834 0 _0102_
rlabel metal2 24150 6494 24150 6494 0 _0103_
rlabel metal1 21666 3162 21666 3162 0 _0104_
rlabel metal1 21075 6698 21075 6698 0 _0105_
rlabel metal2 20470 3298 20470 3298 0 _0106_
rlabel metal1 19182 3502 19182 3502 0 _0107_
rlabel metal2 13846 2856 13846 2856 0 _0108_
rlabel metal2 14214 6120 14214 6120 0 _0109_
rlabel metal2 13018 3672 13018 3672 0 _0110_
rlabel metal1 17303 3434 17303 3434 0 _0111_
rlabel metal1 17756 6426 17756 6426 0 _0112_
rlabel metal1 18131 3094 18131 3094 0 _0113_
rlabel metal1 15824 10438 15824 10438 0 _0114_
rlabel metal1 15732 15334 15732 15334 0 _0115_
rlabel metal1 16061 11798 16061 11798 0 _0116_
rlabel metal2 15410 13090 15410 13090 0 _0117_
rlabel metal1 18216 15674 18216 15674 0 _0118_
rlabel metal1 17848 11322 17848 11322 0 _0119_
rlabel metal2 20102 14552 20102 14552 0 _0120_
rlabel metal2 20286 14382 20286 14382 0 _0121_
rlabel metal1 20976 15130 20976 15130 0 _0122_
rlabel metal1 17664 16558 17664 16558 0 _0123_
rlabel metal2 22770 17000 22770 17000 0 _0124_
rlabel metal1 23506 17136 23506 17136 0 _0125_
rlabel metal1 23835 18666 23835 18666 0 _0126_
rlabel metal1 23276 19482 23276 19482 0 _0127_
rlabel metal1 21351 20842 21351 20842 0 _0128_
rlabel metal1 23644 25466 23644 25466 0 _0129_
rlabel metal1 24012 20774 24012 20774 0 _0130_
rlabel metal2 23782 22372 23782 22372 0 _0131_
rlabel metal1 24479 23766 24479 23766 0 _0132_
rlabel metal1 21397 22678 21397 22678 0 _0133_
rlabel metal1 20700 26282 20700 26282 0 _0134_
rlabel metal1 20516 26418 20516 26418 0 _0135_
rlabel metal2 13846 26180 13846 26180 0 _0136_
rlabel metal2 14398 21352 14398 21352 0 _0137_
rlabel metal1 13064 23834 13064 23834 0 _0138_
rlabel metal2 12742 25704 12742 25704 0 _0139_
rlabel metal1 15456 26282 15456 26282 0 _0140_
rlabel metal1 18775 25942 18775 25942 0 _0141_
rlabel metal2 19182 24990 19182 24990 0 _0142_
rlabel metal2 11638 25466 11638 25466 0 _0143_
rlabel metal2 13110 21522 13110 21522 0 _0144_
rlabel metal2 7498 25874 7498 25874 0 _0145_
rlabel metal2 6946 25704 6946 25704 0 _0146_
rlabel metal2 11638 24004 11638 24004 0 _0147_
rlabel metal1 5980 24786 5980 24786 0 _0148_
rlabel metal2 6578 23970 6578 23970 0 _0149_
rlabel metal2 5198 18122 5198 18122 0 _0150_
rlabel metal1 9706 19754 9706 19754 0 _0151_
rlabel metal1 9798 19278 9798 19278 0 _0152_
rlabel metal1 6532 14586 6532 14586 0 _0153_
rlabel metal2 4094 22882 4094 22882 0 _0154_
rlabel metal1 9246 14314 9246 14314 0 _0155_
rlabel metal1 7774 16218 7774 16218 0 _0156_
rlabel metal1 4876 16762 4876 16762 0 _0157_
rlabel metal1 8464 19482 8464 19482 0 _0158_
rlabel metal1 8464 17102 8464 17102 0 _0159_
rlabel metal2 8970 21726 8970 21726 0 _0160_
rlabel metal1 8602 21896 8602 21896 0 _0161_
rlabel metal1 9660 15062 9660 15062 0 _0162_
rlabel metal2 7406 14178 7406 14178 0 _0163_
rlabel metal2 1702 15470 1702 15470 0 _0164_
rlabel metal1 2070 15538 2070 15538 0 _0165_
rlabel metal2 4922 14756 4922 14756 0 _0166_
rlabel metal2 1702 17816 1702 17816 0 _0167_
rlabel metal2 2162 21284 2162 21284 0 _0168_
rlabel metal2 1702 19550 1702 19550 0 _0169_
rlabel metal2 5934 20434 5934 20434 0 _0170_
rlabel metal2 6670 21726 6670 21726 0 _0171_
rlabel metal1 3864 21114 3864 21114 0 _0172_
rlabel metal1 8500 9554 8500 9554 0 _0173_
rlabel metal1 11270 6290 11270 6290 0 _0174_
rlabel metal1 10150 3094 10150 3094 0 _0175_
rlabel metal1 10897 3502 10897 3502 0 _0176_
rlabel metal2 12742 6562 12742 6562 0 _0177_
rlabel metal2 8970 6902 8970 6902 0 _0178_
rlabel metal1 3864 17578 3864 17578 0 _0179_
rlabel via1 8413 4114 8413 4114 0 _0180_
rlabel metal1 8648 3162 8648 3162 0 _0181_
rlabel metal1 5975 3434 5975 3434 0 _0182_
rlabel metal1 4912 3026 4912 3026 0 _0183_
rlabel via1 4641 4182 4641 4182 0 _0184_
rlabel via1 10161 8874 10161 8874 0 _0185_
rlabel metal1 7866 11798 7866 11798 0 _0186_
rlabel metal2 2530 11866 2530 11866 0 _0187_
rlabel metal1 2208 11594 2208 11594 0 _0188_
rlabel metal1 5750 13362 5750 13362 0 _0189_
rlabel metal1 4273 12818 4273 12818 0 _0190_
rlabel metal1 8188 8058 8188 8058 0 _0191_
rlabel metal1 7125 9554 7125 9554 0 _0192_
rlabel metal1 4411 6698 4411 6698 0 _0193_
rlabel metal1 2346 7480 2346 7480 0 _0194_
rlabel metal1 2208 9146 2208 9146 0 _0195_
rlabel metal1 2238 9962 2238 9962 0 _0196_
rlabel metal1 8091 11050 8091 11050 0 _0197_
rlabel metal1 5980 13702 5980 13702 0 _0198_
rlabel metal1 6118 13804 6118 13804 0 _0199_
rlabel metal2 7682 7412 7682 7412 0 _0200_
rlabel metal2 5106 8942 5106 8942 0 _0201_
rlabel viali 5014 8943 5014 8943 0 _0202_
rlabel metal1 5520 9010 5520 9010 0 _0203_
rlabel metal1 7636 10030 7636 10030 0 _0204_
rlabel metal1 4600 7242 4600 7242 0 _0205_
rlabel metal1 4784 7378 4784 7378 0 _0206_
rlabel metal2 1886 9248 1886 9248 0 _0207_
rlabel metal1 3450 7990 3450 7990 0 _0208_
rlabel metal1 3320 7718 3320 7718 0 _0209_
rlabel metal2 3634 7548 3634 7548 0 _0210_
rlabel via1 2538 8874 2538 8874 0 _0211_
rlabel metal1 2484 8942 2484 8942 0 _0212_
rlabel metal2 2898 9928 2898 9928 0 _0213_
rlabel metal2 2806 10234 2806 10234 0 _0214_
rlabel metal1 9016 20910 9016 20910 0 _0215_
rlabel metal1 4646 19822 4646 19822 0 _0216_
rlabel metal2 4462 18700 4462 18700 0 _0217_
rlabel metal1 3864 18258 3864 18258 0 _0218_
rlabel metal2 5934 21556 5934 21556 0 _0219_
rlabel metal1 5612 17646 5612 17646 0 _0220_
rlabel metal1 6540 17238 6540 17238 0 _0221_
rlabel metal2 5750 21182 5750 21182 0 _0222_
rlabel metal2 7498 21250 7498 21250 0 _0223_
rlabel metal1 6026 22032 6026 22032 0 _0224_
rlabel metal1 5750 20434 5750 20434 0 _0225_
rlabel metal2 6118 20026 6118 20026 0 _0226_
rlabel metal2 3450 19482 3450 19482 0 _0227_
rlabel metal1 2714 21046 2714 21046 0 _0228_
rlabel metal1 2622 19754 2622 19754 0 _0229_
rlabel metal1 2438 19856 2438 19856 0 _0230_
rlabel metal1 3450 18190 3450 18190 0 _0231_
rlabel metal1 2484 18258 2484 18258 0 _0232_
rlabel metal1 5842 18224 5842 18224 0 _0233_
rlabel metal1 5566 16048 5566 16048 0 _0234_
rlabel metal1 5152 14382 5152 14382 0 _0235_
rlabel metal2 4002 16218 4002 16218 0 _0236_
rlabel metal1 2898 16116 2898 16116 0 _0237_
rlabel metal1 5474 20570 5474 20570 0 _0238_
rlabel metal1 4508 15538 4508 15538 0 _0239_
rlabel metal2 2346 15878 2346 15878 0 _0240_
rlabel metal2 17894 7548 17894 7548 0 _0241_
rlabel metal1 16974 10166 16974 10166 0 _0242_
rlabel metal1 7544 15538 7544 15538 0 _0243_
rlabel metal1 7452 13906 7452 13906 0 _0244_
rlabel metal1 14674 11322 14674 11322 0 _0245_
rlabel metal2 8970 15946 8970 15946 0 _0246_
rlabel metal1 9154 14790 9154 14790 0 _0247_
rlabel metal1 15088 21386 15088 21386 0 _0248_
rlabel metal1 8878 21114 8878 21114 0 _0249_
rlabel metal1 13432 21862 13432 21862 0 _0250_
rlabel metal2 8050 21250 8050 21250 0 _0251_
rlabel metal1 8786 21658 8786 21658 0 _0252_
rlabel metal2 8786 18394 8786 18394 0 _0253_
rlabel metal1 9246 18190 9246 18190 0 _0254_
rlabel metal1 8602 19924 8602 19924 0 _0255_
rlabel metal1 8326 19346 8326 19346 0 _0256_
rlabel metal1 6118 16626 6118 16626 0 _0257_
rlabel metal1 5244 16558 5244 16558 0 _0258_
rlabel metal1 6900 17578 6900 17578 0 _0259_
rlabel metal1 7452 17714 7452 17714 0 _0260_
rlabel metal2 8418 16932 8418 16932 0 _0261_
rlabel metal1 12558 9520 12558 9520 0 _0262_
rlabel metal1 9062 13804 9062 13804 0 _0263_
rlabel metal1 8832 14042 8832 14042 0 _0264_
rlabel metal1 5198 22508 5198 22508 0 _0265_
rlabel metal1 4416 22610 4416 22610 0 _0266_
rlabel metal1 6946 15980 6946 15980 0 _0267_
rlabel metal1 6486 14382 6486 14382 0 _0268_
rlabel metal2 10350 19091 10350 19091 0 _0269_
rlabel metal1 9752 18938 9752 18938 0 _0270_
rlabel metal1 4738 20026 4738 20026 0 _0271_
rlabel metal1 10718 20332 10718 20332 0 _0272_
rlabel metal2 9614 20060 9614 20060 0 _0273_
rlabel metal2 21574 11373 21574 11373 0 _0274_
rlabel metal1 21758 11085 21758 11085 0 _0275_
rlabel metal1 21298 10982 21298 10982 0 _0276_
rlabel metal1 23246 9962 23246 9962 0 _0277_
rlabel metal1 21130 11050 21130 11050 0 _0278_
rlabel metal2 22034 11084 22034 11084 0 _0279_
rlabel metal1 23966 10132 23966 10132 0 _0280_
rlabel metal1 23966 11084 23966 11084 0 _0281_
rlabel metal1 23782 11118 23782 11118 0 _0282_
rlabel metal1 24380 10234 24380 10234 0 _0283_
rlabel metal1 24886 10234 24886 10234 0 _0284_
rlabel metal1 24748 10710 24748 10710 0 _0285_
rlabel metal2 21390 9724 21390 9724 0 _0286_
rlabel metal2 21482 10064 21482 10064 0 _0287_
rlabel metal1 22356 11186 22356 11186 0 _0288_
rlabel metal2 22310 9996 22310 9996 0 _0289_
rlabel metal1 21574 10710 21574 10710 0 _0290_
rlabel metal2 21206 11492 21206 11492 0 _0291_
rlabel metal1 21666 11730 21666 11730 0 _0292_
rlabel metal1 21574 11628 21574 11628 0 _0293_
rlabel metal1 21712 11866 21712 11866 0 _0294_
rlabel metal2 20010 6222 20010 6222 0 _0295_
rlabel metal1 21022 4624 21022 4624 0 _0296_
rlabel metal1 20516 4658 20516 4658 0 _0297_
rlabel metal1 21988 5610 21988 5610 0 _0298_
rlabel metal2 19458 3740 19458 3740 0 _0299_
rlabel metal1 20746 5338 20746 5338 0 _0300_
rlabel metal1 22218 5678 22218 5678 0 _0301_
rlabel metal1 22632 5882 22632 5882 0 _0302_
rlabel metal2 22678 5678 22678 5678 0 _0303_
rlabel metal1 22816 4046 22816 4046 0 _0304_
rlabel metal1 22126 4624 22126 4624 0 _0305_
rlabel metal1 22678 4182 22678 4182 0 _0306_
rlabel metal2 19274 6460 19274 6460 0 _0307_
rlabel metal1 20562 6256 20562 6256 0 _0308_
rlabel metal1 20562 5882 20562 5882 0 _0309_
rlabel metal2 21298 6732 21298 6732 0 _0310_
rlabel metal1 20608 6358 20608 6358 0 _0311_
rlabel metal1 19412 5270 19412 5270 0 _0312_
rlabel metal1 20240 4046 20240 4046 0 _0313_
rlabel metal2 20286 3638 20286 3638 0 _0314_
rlabel metal1 20746 4012 20746 4012 0 _0315_
rlabel metal1 19826 4590 19826 4590 0 _0316_
rlabel metal1 15686 6120 15686 6120 0 _0317_
rlabel metal1 17304 5202 17304 5202 0 _0318_
rlabel metal1 16652 5338 16652 5338 0 _0319_
rlabel metal1 14352 4998 14352 4998 0 _0320_
rlabel metal1 15364 5202 15364 5202 0 _0321_
rlabel metal1 15226 5746 15226 5746 0 _0322_
rlabel metal1 14490 3910 14490 3910 0 _0323_
rlabel metal1 14398 4658 14398 4658 0 _0324_
rlabel metal1 14674 3502 14674 3502 0 _0325_
rlabel metal1 15594 3536 15594 3536 0 _0326_
rlabel metal1 14674 4046 14674 4046 0 _0327_
rlabel metal2 15410 3978 15410 3978 0 _0328_
rlabel metal1 14996 6290 14996 6290 0 _0329_
rlabel metal1 15548 6426 15548 6426 0 _0330_
rlabel metal2 16422 5440 16422 5440 0 _0331_
rlabel metal1 15502 5712 15502 5712 0 _0332_
rlabel metal1 15318 5882 15318 5882 0 _0333_
rlabel metal1 17480 4182 17480 4182 0 _0334_
rlabel metal2 16882 4284 16882 4284 0 _0335_
rlabel metal1 17342 4012 17342 4012 0 _0336_
rlabel metal1 16330 5134 16330 5134 0 _0337_
rlabel metal1 18078 13362 18078 13362 0 _0338_
rlabel metal2 18354 14076 18354 14076 0 _0339_
rlabel metal1 17526 14450 17526 14450 0 _0340_
rlabel via1 17258 13974 17258 13974 0 _0341_
rlabel metal1 18278 13974 18278 13974 0 _0342_
rlabel metal2 17342 14688 17342 14688 0 _0343_
rlabel metal2 15962 13906 15962 13906 0 _0344_
rlabel metal1 15778 14382 15778 14382 0 _0345_
rlabel metal1 15134 14416 15134 14416 0 _0346_
rlabel metal2 17618 15572 17618 15572 0 _0347_
rlabel metal1 16928 15062 16928 15062 0 _0348_
rlabel metal2 17066 15266 17066 15266 0 _0349_
rlabel metal1 17066 12240 17066 12240 0 _0350_
rlabel metal1 17112 12410 17112 12410 0 _0351_
rlabel metal1 17848 13226 17848 13226 0 _0352_
rlabel metal1 17250 12954 17250 12954 0 _0353_
rlabel metal1 16882 13328 16882 13328 0 _0354_
rlabel metal1 20010 13430 20010 13430 0 _0355_
rlabel metal2 18538 14586 18538 14586 0 _0356_
rlabel metal1 18814 14042 18814 14042 0 _0357_
rlabel metal2 18630 13056 18630 13056 0 _0358_
rlabel via1 20746 19261 20746 19261 0 _0359_
rlabel metal1 21482 19380 21482 19380 0 _0360_
rlabel via1 21587 19754 21587 19754 0 _0361_
rlabel metal1 19734 17068 19734 17068 0 _0362_
rlabel metal1 22218 19346 22218 19346 0 _0363_
rlabel metal1 20792 17578 20792 17578 0 _0364_
rlabel metal2 20562 16830 20562 16830 0 _0365_
rlabel via2 21298 16541 21298 16541 0 _0366_
rlabel metal1 21482 16150 21482 16150 0 _0367_
rlabel metal1 20838 17136 20838 17136 0 _0368_
rlabel metal2 20010 17340 20010 17340 0 _0369_
rlabel metal1 21160 17578 21160 17578 0 _0370_
rlabel metal1 21206 18292 21206 18292 0 _0371_
rlabel metal2 21390 18564 21390 18564 0 _0372_
rlabel metal1 21114 20366 21114 20366 0 _0373_
rlabel metal2 21114 18428 21114 18428 0 _0374_
rlabel metal1 20976 18394 20976 18394 0 _0375_
rlabel metal2 21390 20026 21390 20026 0 _0376_
rlabel metal2 21298 19652 21298 19652 0 _0377_
rlabel metal1 21390 19890 21390 19890 0 _0378_
rlabel metal1 20470 19482 20470 19482 0 _0379_
rlabel via1 20194 23069 20194 23069 0 _0380_
rlabel viali 21574 24789 21574 24789 0 _0381_
rlabel metal1 20976 24582 20976 24582 0 _0382_
rlabel metal1 21935 23018 21935 23018 0 _0383_
rlabel metal1 21298 24174 21298 24174 0 _0384_
rlabel metal1 20746 23664 20746 23664 0 _0385_
rlabel metal1 23736 23154 23736 23154 0 _0386_
rlabel metal1 23276 23290 23276 23290 0 _0387_
rlabel metal2 22218 23970 22218 23970 0 _0388_
rlabel metal1 23690 23290 23690 23290 0 _0389_
rlabel metal1 22632 23290 22632 23290 0 _0390_
rlabel metal2 22954 23970 22954 23970 0 _0391_
rlabel metal2 19734 22916 19734 22916 0 _0392_
rlabel metal1 20654 23120 20654 23120 0 _0393_
rlabel metal1 21068 24242 21068 24242 0 _0394_
rlabel metal1 20976 23290 20976 23290 0 _0395_
rlabel metal2 20470 23290 20470 23290 0 _0396_
rlabel metal1 20930 24378 20930 24378 0 _0397_
rlabel metal2 20562 24548 20562 24548 0 _0398_
rlabel metal1 21022 24820 21022 24820 0 _0399_
rlabel metal1 20194 24684 20194 24684 0 _0400_
rlabel metal1 18170 24616 18170 24616 0 _0401_
rlabel metal2 18262 25228 18262 25228 0 _0402_
rlabel metal1 17460 24888 17460 24888 0 _0403_
rlabel metal1 13938 24242 13938 24242 0 _0404_
rlabel metal1 16698 24752 16698 24752 0 _0405_
rlabel metal1 14904 24786 14904 24786 0 _0406_
rlabel metal2 13938 24208 13938 24208 0 _0407_
rlabel metal2 13846 25092 13846 25092 0 _0408_
rlabel metal1 13248 24854 13248 24854 0 _0409_
rlabel metal1 14352 23562 14352 23562 0 _0410_
rlabel metal2 14674 24582 14674 24582 0 _0411_
rlabel metal1 14306 24752 14306 24752 0 _0412_
rlabel metal1 15180 24378 15180 24378 0 _0413_
rlabel metal1 15410 24922 15410 24922 0 _0414_
rlabel metal2 16790 24956 16790 24956 0 _0415_
rlabel metal1 16008 24378 16008 24378 0 _0416_
rlabel metal1 15134 25296 15134 25296 0 _0417_
rlabel metal1 17526 24310 17526 24310 0 _0418_
rlabel metal2 17802 25585 17802 25585 0 _0419_
rlabel metal1 17342 24718 17342 24718 0 _0420_
rlabel metal2 18446 25602 18446 25602 0 _0421_
rlabel metal1 7544 24786 7544 24786 0 _0422_
rlabel metal2 8970 24140 8970 24140 0 _0423_
rlabel metal1 9890 26316 9890 26316 0 _0424_
rlabel metal1 9108 25194 9108 25194 0 _0425_
rlabel metal2 7866 24276 7866 24276 0 _0426_
rlabel metal2 9430 25976 9430 25976 0 _0427_
rlabel metal2 9614 25534 9614 25534 0 _0428_
rlabel metal1 9890 25466 9890 25466 0 _0429_
rlabel metal1 9798 25262 9798 25262 0 _0430_
rlabel metal1 10442 25738 10442 25738 0 _0431_
rlabel metal1 9154 25806 9154 25806 0 _0432_
rlabel metal1 9476 25942 9476 25942 0 _0433_
rlabel metal1 9706 23086 9706 23086 0 _0434_
rlabel metal2 9890 23732 9890 23732 0 _0435_
rlabel metal2 8510 24140 8510 24140 0 _0436_
rlabel metal1 9936 23834 9936 23834 0 _0437_
rlabel metal1 9338 24106 9338 24106 0 _0438_
rlabel metal1 8050 23834 8050 23834 0 _0439_
rlabel metal1 7828 24184 7828 24184 0 _0440_
rlabel metal2 8188 24174 8188 24174 0 _0441_
rlabel metal2 7314 24140 7314 24140 0 _0442_
rlabel metal1 5060 23698 5060 23698 0 _0443_
rlabel metal2 14582 17612 14582 17612 0 _0444_
rlabel metal2 13662 19924 13662 19924 0 _0445_
rlabel metal1 13018 20400 13018 20400 0 _0446_
rlabel metal2 14030 19618 14030 19618 0 _0447_
rlabel metal1 14122 14280 14122 14280 0 _0448_
rlabel metal1 10626 12784 10626 12784 0 _0449_
rlabel via2 14490 18853 14490 18853 0 _0450_
rlabel metal1 13846 17850 13846 17850 0 _0451_
rlabel metal1 14536 17646 14536 17646 0 _0452_
rlabel metal1 11546 13226 11546 13226 0 _0453_
rlabel metal1 14858 17136 14858 17136 0 _0454_
rlabel metal2 14490 15028 14490 15028 0 _0455_
rlabel metal1 12934 17510 12934 17510 0 _0456_
rlabel metal2 13478 16422 13478 16422 0 _0457_
rlabel metal1 11546 18326 11546 18326 0 _0458_
rlabel metal2 10350 16354 10350 16354 0 _0459_
rlabel metal1 9982 16558 9982 16558 0 _0460_
rlabel metal1 11914 16626 11914 16626 0 _0461_
rlabel metal1 10304 17306 10304 17306 0 _0462_
rlabel metal2 12742 16660 12742 16660 0 _0463_
rlabel metal2 11546 17442 11546 17442 0 _0464_
rlabel metal2 11454 17068 11454 17068 0 _0465_
rlabel metal1 13110 17816 13110 17816 0 _0466_
rlabel metal1 13248 17850 13248 17850 0 _0467_
rlabel metal1 12006 18156 12006 18156 0 _0468_
rlabel metal1 11408 18190 11408 18190 0 _0469_
rlabel metal1 10580 16082 10580 16082 0 _0470_
rlabel metal1 11040 16218 11040 16218 0 _0471_
rlabel metal2 12466 10370 12466 10370 0 _0472_
rlabel metal1 9660 12750 9660 12750 0 _0473_
rlabel metal1 12006 13294 12006 13294 0 _0474_
rlabel metal1 10672 13906 10672 13906 0 _0475_
rlabel metal1 11362 14042 11362 14042 0 _0476_
rlabel metal2 12374 13804 12374 13804 0 _0477_
rlabel metal1 12604 13498 12604 13498 0 _0478_
rlabel metal2 11914 15300 11914 15300 0 _0479_
rlabel metal2 12558 14790 12558 14790 0 _0480_
rlabel metal1 23322 17646 23322 17646 0 _0481_
rlabel metal2 13294 19516 13294 19516 0 _0482_
rlabel metal1 12788 19822 12788 19822 0 _0483_
rlabel metal2 9154 20213 9154 20213 0 _0484_
rlabel metal2 2346 19822 2346 19822 0 _0485_
rlabel metal2 5198 10268 5198 10268 0 _0486_
rlabel metal2 1794 9316 1794 9316 0 _0487_
rlabel metal1 6210 9044 6210 9044 0 _0488_
rlabel metal2 6302 8296 6302 8296 0 _0489_
rlabel metal1 5842 8432 5842 8432 0 _0490_
rlabel metal1 5842 7922 5842 7922 0 _0491_
rlabel metal1 5152 8602 5152 8602 0 _0492_
rlabel metal1 6210 8942 6210 8942 0 _0493_
rlabel metal2 5566 9690 5566 9690 0 _0494_
rlabel metal1 4462 9146 4462 9146 0 _0495_
rlabel metal1 5428 9486 5428 9486 0 _0496_
rlabel metal2 6394 9418 6394 9418 0 _0497_
rlabel metal1 18262 21114 18262 21114 0 _0498_
rlabel metal1 18492 22610 18492 22610 0 _0499_
rlabel metal1 17434 21930 17434 21930 0 _0500_
rlabel metal1 18078 22678 18078 22678 0 _0501_
rlabel metal1 18538 22542 18538 22542 0 _0502_
rlabel metal2 17756 21828 17756 21828 0 _0503_
rlabel metal2 18078 19788 18078 19788 0 _0504_
rlabel metal2 25162 19380 25162 19380 0 _0505_
rlabel metal1 17664 22474 17664 22474 0 _0506_
rlabel metal2 18998 21726 18998 21726 0 _0507_
rlabel metal1 18216 21386 18216 21386 0 _0508_
rlabel metal1 18308 21522 18308 21522 0 _0509_
rlabel metal2 17894 20570 17894 20570 0 _0510_
rlabel metal1 17020 19210 17020 19210 0 _0511_
rlabel metal1 17710 18734 17710 18734 0 _0512_
rlabel metal1 17618 19482 17618 19482 0 _0513_
rlabel metal2 17250 19210 17250 19210 0 _0514_
rlabel metal1 2507 17238 2507 17238 0 _0515_
rlabel metal2 15962 22610 15962 22610 0 _0516_
rlabel metal1 15410 22066 15410 22066 0 _0517_
rlabel metal1 15870 21930 15870 21930 0 _0518_
rlabel metal1 16192 21862 16192 21862 0 _0519_
rlabel metal1 17986 18258 17986 18258 0 _0520_
rlabel metal2 16514 18496 16514 18496 0 _0521_
rlabel metal1 17158 3162 17158 3162 0 _0522_
rlabel metal1 17434 22202 17434 22202 0 _0523_
rlabel metal1 16238 22134 16238 22134 0 _0524_
rlabel metal1 17204 17646 17204 17646 0 _0525_
rlabel metal1 18367 18394 18367 18394 0 _0526_
rlabel metal1 17158 18054 17158 18054 0 _0527_
rlabel metal2 16882 18428 16882 18428 0 _0528_
rlabel metal1 16974 17850 16974 17850 0 _0529_
rlabel metal1 15962 18598 15962 18598 0 _0530_
rlabel metal1 17158 20502 17158 20502 0 _0531_
rlabel metal1 17434 21658 17434 21658 0 _0532_
rlabel metal1 16238 22066 16238 22066 0 _0533_
rlabel metal2 16238 22474 16238 22474 0 _0534_
rlabel metal1 16806 20842 16806 20842 0 _0535_
rlabel metal1 16054 20842 16054 20842 0 _0536_
rlabel metal1 16698 19890 16698 19890 0 _0537_
rlabel metal2 16054 20774 16054 20774 0 _0538_
rlabel metal2 16330 20026 16330 20026 0 _0539_
rlabel metal2 16514 20077 16514 20077 0 _0540_
rlabel metal1 16192 18734 16192 18734 0 _0541_
rlabel metal1 16330 18394 16330 18394 0 _0542_
rlabel metal1 17250 18768 17250 18768 0 _0543_
rlabel metal1 13662 15096 13662 15096 0 _0544_
rlabel metal2 2346 8636 2346 8636 0 _0545_
rlabel metal1 16100 19346 16100 19346 0 _0546_
rlabel metal1 16238 19176 16238 19176 0 _0547_
rlabel metal2 12834 14246 12834 14246 0 _0548_
rlabel metal2 2714 11951 2714 11951 0 _0549_
rlabel metal1 7544 9146 7544 9146 0 _0550_
rlabel metal1 23874 12818 23874 12818 0 _0551_
rlabel metal1 21252 3026 21252 3026 0 _0552_
rlabel metal1 15456 12818 15456 12818 0 _0553_
rlabel metal1 24012 21998 24012 21998 0 _0554_
rlabel metal2 19458 20383 19458 20383 0 _0555_
rlabel metal1 14904 18054 14904 18054 0 _0556_
rlabel metal1 16192 10234 16192 10234 0 _0557_
rlabel metal1 19504 10438 19504 10438 0 _0558_
rlabel metal1 18216 10166 18216 10166 0 _0559_
rlabel metal2 18446 10812 18446 10812 0 _0560_
rlabel metal1 18538 10608 18538 10608 0 _0561_
rlabel metal1 14858 11152 14858 11152 0 _0562_
rlabel via1 14398 10642 14398 10642 0 _0563_
rlabel metal1 13478 10064 13478 10064 0 _0564_
rlabel metal2 13984 17612 13984 17612 0 _0565_
rlabel metal2 19458 11322 19458 11322 0 _0566_
rlabel metal1 18998 9588 18998 9588 0 _0567_
rlabel metal1 16698 9690 16698 9690 0 _0568_
rlabel metal1 19274 9520 19274 9520 0 _0569_
rlabel metal2 18722 10336 18722 10336 0 _0570_
rlabel metal1 14214 11186 14214 11186 0 _0571_
rlabel metal1 14582 10234 14582 10234 0 _0572_
rlabel metal1 12788 10030 12788 10030 0 _0573_
rlabel metal1 15640 9350 15640 9350 0 _0574_
rlabel metal2 16330 9044 16330 9044 0 _0575_
rlabel metal1 15962 9622 15962 9622 0 _0576_
rlabel metal1 12926 10064 12926 10064 0 _0577_
rlabel metal2 12650 9486 12650 9486 0 _0578_
rlabel metal1 13386 9486 13386 9486 0 _0579_
rlabel metal1 15916 8058 15916 8058 0 _0580_
rlabel metal2 18078 8194 18078 8194 0 _0581_
rlabel metal2 16698 8840 16698 8840 0 _0582_
rlabel metal1 13570 7820 13570 7820 0 _0583_
rlabel metal1 13754 7990 13754 7990 0 _0584_
rlabel metal1 12834 7854 12834 7854 0 _0585_
rlabel metal2 12926 8806 12926 8806 0 _0586_
rlabel via1 13202 9622 13202 9622 0 _0587_
rlabel metal1 14030 9622 14030 9622 0 _0588_
rlabel metal1 13938 8874 13938 8874 0 _0589_
rlabel metal1 18400 8466 18400 8466 0 _0590_
rlabel metal1 18492 7514 18492 7514 0 _0591_
rlabel metal2 19182 7922 19182 7922 0 _0592_
rlabel metal2 18170 8636 18170 8636 0 _0593_
rlabel metal1 15456 9146 15456 9146 0 _0594_
rlabel metal1 13156 8874 13156 8874 0 _0595_
rlabel metal1 17940 9146 17940 9146 0 _0596_
rlabel metal1 18492 7990 18492 7990 0 _0597_
rlabel metal2 19734 8568 19734 8568 0 _0598_
rlabel metal2 18078 9418 18078 9418 0 _0599_
rlabel metal1 13018 8874 13018 8874 0 _0600_
rlabel metal1 13570 8500 13570 8500 0 _0601_
rlabel metal1 13432 9146 13432 9146 0 _0602_
rlabel metal2 14122 9350 14122 9350 0 _0603_
rlabel metal1 13754 9690 13754 9690 0 _0604_
rlabel metal1 13616 10642 13616 10642 0 _0605_
rlabel metal2 13202 10234 13202 10234 0 _0606_
rlabel metal2 12742 8670 12742 8670 0 _0607_
rlabel metal2 13938 8262 13938 8262 0 _0608_
rlabel metal1 13662 9418 13662 9418 0 _0609_
rlabel metal1 14260 8262 14260 8262 0 _0610_
rlabel metal1 12558 8296 12558 8296 0 _0611_
rlabel metal1 9798 7310 9798 7310 0 _0612_
rlabel metal1 10304 6222 10304 6222 0 _0613_
rlabel metal1 10902 5134 10902 5134 0 _0614_
rlabel metal1 9108 5610 9108 5610 0 _0615_
rlabel viali 9246 5678 9246 5678 0 _0616_
rlabel metal1 8970 5678 8970 5678 0 _0617_
rlabel metal1 9890 5882 9890 5882 0 _0618_
rlabel metal2 10074 6018 10074 6018 0 _0619_
rlabel metal1 9568 6290 9568 6290 0 _0620_
rlabel metal1 10304 6426 10304 6426 0 _0621_
rlabel metal1 10902 6970 10902 6970 0 _0622_
rlabel metal1 10166 7854 10166 7854 0 _0623_
rlabel metal1 10626 6834 10626 6834 0 _0624_
rlabel metal1 10028 7718 10028 7718 0 _0625_
rlabel metal1 9982 7922 9982 7922 0 _0626_
rlabel metal2 10994 4896 10994 4896 0 _0627_
rlabel metal2 11914 4454 11914 4454 0 _0628_
rlabel metal2 10074 4352 10074 4352 0 _0629_
rlabel metal1 11086 3978 11086 3978 0 _0630_
rlabel metal2 11362 5950 11362 5950 0 _0631_
rlabel metal1 10948 5338 10948 5338 0 _0632_
rlabel metal1 7130 4998 7130 4998 0 _0633_
rlabel metal2 6578 4250 6578 4250 0 _0634_
rlabel metal2 7682 6052 7682 6052 0 _0635_
rlabel metal2 6578 6460 6578 6460 0 _0636_
rlabel metal2 7590 5950 7590 5950 0 _0637_
rlabel metal1 7314 6290 7314 6290 0 _0638_
rlabel metal1 5842 6392 5842 6392 0 _0639_
rlabel metal2 6946 5916 6946 5916 0 _0640_
rlabel metal1 6072 5338 6072 5338 0 _0641_
rlabel metal1 5566 6256 5566 6256 0 _0642_
rlabel via1 7230 5338 7230 5338 0 _0643_
rlabel metal1 7912 4590 7912 4590 0 _0644_
rlabel metal2 7866 6154 7866 6154 0 _0645_
rlabel metal2 7682 5066 7682 5066 0 _0646_
rlabel metal1 7828 4250 7828 4250 0 _0647_
rlabel metal1 8280 3910 8280 3910 0 _0648_
rlabel metal1 8472 3434 8472 3434 0 _0649_
rlabel metal2 8694 3332 8694 3332 0 _0650_
rlabel metal1 5842 4590 5842 4590 0 _0651_
rlabel metal2 6670 3400 6670 3400 0 _0652_
rlabel metal1 6808 3162 6808 3162 0 _0653_
rlabel metal2 6210 3162 6210 3162 0 _0654_
rlabel metal1 6448 3366 6448 3366 0 _0655_
rlabel via2 4922 3485 4922 3485 0 _0656_
rlabel metal1 6080 4454 6080 4454 0 _0657_
rlabel metal1 5198 4624 5198 4624 0 _0658_
rlabel metal1 7084 13498 7084 13498 0 _0659_
rlabel metal2 4830 12648 4830 12648 0 _0660_
rlabel metal2 3910 11900 3910 11900 0 _0661_
rlabel metal2 6026 11492 6026 11492 0 _0662_
rlabel metal1 6440 11322 6440 11322 0 _0663_
rlabel metal2 4922 11526 4922 11526 0 _0664_
rlabel metal2 5842 12002 5842 12002 0 _0665_
rlabel metal1 6256 11866 6256 11866 0 _0666_
rlabel metal2 5474 11764 5474 11764 0 _0667_
rlabel metal1 7460 13158 7460 13158 0 _0668_
rlabel metal1 6394 13328 6394 13328 0 _0669_
rlabel metal2 7406 13260 7406 13260 0 _0670_
rlabel metal1 7314 12614 7314 12614 0 _0671_
rlabel metal1 4278 11322 4278 11322 0 _0672_
rlabel metal1 2898 11696 2898 11696 0 _0673_
rlabel metal1 2760 11798 2760 11798 0 _0674_
rlabel metal1 2116 11798 2116 11798 0 _0675_
rlabel metal2 5290 18530 5290 18530 0 clknet_0_CLK_SR
rlabel metal2 19090 18292 19090 18292 0 clknet_0_Dead_Time_Generator_inst_1.clk
rlabel metal1 1426 17680 1426 17680 0 clknet_1_0__leaf_CLK_SR
rlabel metal1 1472 21454 1472 21454 0 clknet_1_1__leaf_CLK_SR
rlabel metal1 2622 7242 2622 7242 0 clknet_3_0__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal2 2162 12512 2162 12512 0 clknet_3_1__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal2 21942 6800 21942 6800 0 clknet_3_2__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 14214 11730 14214 11730 0 clknet_3_3__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal2 12098 21760 12098 21760 0 clknet_3_4__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 12006 24174 12006 24174 0 clknet_3_5__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal2 22126 17952 22126 17952 0 clknet_3_6__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal1 22954 20468 22954 20468 0 clknet_3_7__leaf_Dead_Time_Generator_inst_1.clk
rlabel metal2 3910 1588 3910 1588 0 d1[0]
rlabel metal2 7774 1588 7774 1588 0 d1[1]
rlabel metal2 25806 4369 25806 4369 0 d1[2]
rlabel metal2 11638 1588 11638 1588 0 d1[3]
rlabel metal2 25806 21335 25806 21335 0 d1[4]
rlabel via2 25806 25245 25806 25245 0 d1[5]
rlabel metal3 820 21148 820 21148 0 d2[0]
rlabel metal1 15640 26962 15640 26962 0 d2[1]
rlabel metal2 15502 1588 15502 1588 0 d2[2]
rlabel metal3 820 16388 820 16388 0 d2[3]
rlabel metal3 1050 29308 1050 29308 0 d2[4]
rlabel metal2 25806 13141 25806 13141 0 d2[5]
rlabel metal2 1978 11458 1978 11458 0 net1
rlabel metal2 16330 26316 16330 26316 0 net10
rlabel metal1 15962 2618 15962 2618 0 net11
rlabel metal1 1794 16762 1794 16762 0 net12
rlabel metal1 2116 26758 2116 26758 0 net13
rlabel metal1 25530 13498 25530 13498 0 net14
rlabel metal2 14766 17408 14766 17408 0 net15
rlabel metal2 11730 19142 11730 19142 0 net16
rlabel metal1 15088 16966 15088 16966 0 net17
rlabel metal2 23414 26486 23414 26486 0 net18
rlabel metal1 20194 2448 20194 2448 0 net19
rlabel metal1 23782 2618 23782 2618 0 net2
rlabel metal2 25714 16966 25714 16966 0 net20
rlabel metal1 14352 18394 14352 18394 0 net21
rlabel metal1 19550 2346 19550 2346 0 net22
rlabel metal1 1518 12920 1518 12920 0 net23
rlabel metal2 10074 18632 10074 18632 0 net24
rlabel metal1 1518 2448 1518 2448 0 net25
rlabel metal1 7544 2278 7544 2278 0 net3
rlabel metal2 9338 14620 9338 14620 0 net30
rlabel metal1 10212 14042 10212 14042 0 net31
rlabel metal2 9614 11900 9614 11900 0 net32
rlabel metal1 12558 9010 12558 9010 0 net33
rlabel metal1 11592 12410 11592 12410 0 net34
rlabel metal1 9660 11866 9660 11866 0 net35
rlabel metal2 12006 10744 12006 10744 0 net36
rlabel metal1 5382 13974 5382 13974 0 net37
rlabel metal1 8326 12818 8326 12818 0 net38
rlabel via1 10235 6290 10235 6290 0 net39
rlabel metal1 8602 2618 8602 2618 0 net4
rlabel metal1 10350 7378 10350 7378 0 net40
rlabel metal1 14582 18768 14582 18768 0 net41
rlabel metal2 12190 6562 12190 6562 0 net42
rlabel metal1 7866 12682 7866 12682 0 net43
rlabel metal1 8556 12614 8556 12614 0 net44
rlabel metal2 7038 11137 7038 11137 0 net45
rlabel metal1 4812 9554 4812 9554 0 net46
rlabel metal2 6026 9792 6026 9792 0 net47
rlabel metal1 15042 12240 15042 12240 0 net48
rlabel via1 12742 22073 12742 22073 0 net49
rlabel metal1 11638 8942 11638 8942 0 net5
rlabel metal1 9614 6154 9614 6154 0 net50
rlabel metal1 23322 20876 23322 20876 0 net51
rlabel metal2 20286 8772 20286 8772 0 net52
rlabel metal2 5382 8296 5382 8296 0 net53
rlabel metal1 10672 6290 10672 6290 0 net54
rlabel metal2 13202 6120 13202 6120 0 net55
rlabel via2 4738 11747 4738 11747 0 net56
rlabel metal1 15180 21998 15180 21998 0 net57
rlabel metal1 16330 17238 16330 17238 0 net58
rlabel metal1 13662 6732 13662 6732 0 net59
rlabel metal1 12006 2618 12006 2618 0 net6
rlabel metal2 21482 7548 21482 7548 0 net60
rlabel metal2 4002 21114 4002 21114 0 net61
rlabel metal2 14950 24956 14950 24956 0 net62
rlabel metal2 20194 5967 20194 5967 0 net63
rlabel metal1 4048 19890 4048 19890 0 net64
rlabel via2 23138 24157 23138 24157 0 net65
rlabel metal1 15226 3434 15226 3434 0 net66
rlabel metal1 1886 20876 1886 20876 0 net67
rlabel metal2 17250 15028 17250 15028 0 net68
rlabel metal1 21344 19754 21344 19754 0 net69
rlabel metal2 25990 20672 25990 20672 0 net7
rlabel metal2 12650 4352 12650 4352 0 net70
rlabel metal1 5750 12614 5750 12614 0 net71
rlabel metal1 5009 13226 5009 13226 0 net72
rlabel metal1 22080 12818 22080 12818 0 net73
rlabel metal2 3818 11900 3818 11900 0 net74
rlabel metal1 24426 11152 24426 11152 0 net75
rlabel metal1 5658 22746 5658 22746 0 net76
rlabel metal1 18722 14416 18722 14416 0 net77
rlabel metal1 19872 13498 19872 13498 0 net78
rlabel metal1 7452 16082 7452 16082 0 net79
rlabel via2 14674 18275 14674 18275 0 net8
rlabel metal2 21298 18020 21298 18020 0 net80
rlabel metal2 20746 24905 20746 24905 0 net81
rlabel metal1 17066 4080 17066 4080 0 net82
rlabel metal1 16836 26418 16836 26418 0 net83
rlabel metal1 11960 12274 11960 12274 0 net84
rlabel metal2 11546 12988 11546 12988 0 net85
rlabel metal1 4876 13974 4876 13974 0 net86
rlabel metal2 1610 20621 1610 20621 0 net9
<< properties >>
string FIXED_BBOX 0 0 27481 29625
<< end >>
