magic
tech sky130A
magscale 1 2
timestamp 1697513890
<< obsli1 >>
rect 1104 2159 26312 27217
<< obsm1 >>
rect 14 2128 26312 27248
<< metal2 >>
rect 3238 28825 3294 29625
rect 7102 28825 7158 29625
rect 11610 28825 11666 29625
rect 15474 28825 15530 29625
rect 19338 28825 19394 29625
rect 23202 28825 23258 29625
rect 27066 28825 27122 29625
rect 18 0 74 800
rect 3882 0 3938 800
rect 7746 0 7802 800
rect 11610 0 11666 800
rect 15474 0 15530 800
rect 19982 0 20038 800
rect 23846 0 23902 800
<< obsm2 >>
rect 20 28769 3182 29345
rect 3350 28769 7046 29345
rect 7214 28769 11554 29345
rect 11722 28769 15418 29345
rect 15586 28769 19282 29345
rect 19450 28769 23146 29345
rect 23314 28769 27010 29345
rect 20 856 27122 28769
rect 130 31 3826 856
rect 3994 31 7690 856
rect 7858 31 11554 856
rect 11722 31 15418 856
rect 15586 31 19926 856
rect 20094 31 23790 856
rect 23958 31 27122 856
<< metal3 >>
rect 0 29248 800 29368
rect 0 25168 800 25288
rect 26681 25168 27481 25288
rect 0 21088 800 21208
rect 26681 21088 27481 21208
rect 26681 17008 27481 17128
rect 0 16328 800 16448
rect 26681 12928 27481 13048
rect 0 12248 800 12368
rect 0 8168 800 8288
rect 26681 8168 27481 8288
rect 0 4088 800 4208
rect 26681 4088 27481 4208
rect 26681 8 27481 128
<< obsm3 >>
rect 880 29168 27127 29341
rect 800 25368 27127 29168
rect 880 25088 26601 25368
rect 800 21288 27127 25088
rect 880 21008 26601 21288
rect 800 17208 27127 21008
rect 800 16928 26601 17208
rect 800 16528 27127 16928
rect 880 16248 27127 16528
rect 800 13128 27127 16248
rect 800 12848 26601 13128
rect 800 12448 27127 12848
rect 880 12168 27127 12448
rect 800 8368 27127 12168
rect 880 8088 26601 8368
rect 800 4288 27127 8088
rect 880 4008 26601 4288
rect 800 208 27127 4008
rect 800 35 26601 208
<< metal4 >>
rect 4095 2128 4415 27248
rect 4755 2128 5075 27248
rect 10397 2128 10717 27248
rect 11057 2128 11377 27248
rect 16699 2128 17019 27248
rect 17359 2128 17679 27248
rect 23001 2128 23321 27248
rect 23661 2128 23981 27248
<< obsm4 >>
rect 5579 8059 6381 23493
<< metal5 >>
rect 1056 24572 26360 24892
rect 1056 23912 26360 24232
rect 1056 18316 26360 18636
rect 1056 17656 26360 17976
rect 1056 12060 26360 12380
rect 1056 11400 26360 11720
rect 1056 5804 26360 6124
rect 1056 5144 26360 5464
<< labels >>
rlabel metal3 s 0 4088 800 4208 6 CLK_EXT
port 1 nsew
rlabel metal2 s 27066 28825 27122 29625 6 CLK_PLL
port 2 nsew
rlabel metal3 s 0 25168 800 25288 6 CLK_SR
port 3 nsew
rlabel metal3 s 0 8168 800 8288 6 Data_SR
port 4 nsew
rlabel metal2 s 7102 28825 7158 29625 6 NMOS1_PS1
port 5 nsew
rlabel metal2 s 11610 28825 11666 29625 6 NMOS1_PS2
port 6 nsew
rlabel metal3 s 26681 8168 27481 8288 6 NMOS2_PS1
port 7 nsew
rlabel metal2 s 23202 28825 23258 29625 6 NMOS2_PS2
port 8 nsew
rlabel metal2 s 19982 0 20038 800 6 NMOS_PS3
port 9 nsew
rlabel metal3 s 26681 17008 27481 17128 6 PMOS1_PS1
port 10 nsew
rlabel metal2 s 19338 28825 19394 29625 6 PMOS1_PS2
port 11 nsew
rlabel metal3 s 26681 8 27481 128 6 PMOS2_PS1
port 12 nsew
rlabel metal3 s 0 12248 800 12368 6 PMOS2_PS2
port 13 nsew
rlabel metal2 s 3238 28825 3294 29625 6 PMOS_PS3
port 14 nsew
rlabel metal2 s 23846 0 23902 800 6 RST
port 15 nsew
rlabel metal2 s 18 0 74 800 6 SIGNAL_OUTPUT
port 16 nsew
rlabel metal5 s 1056 24572 26360 24892 6 VGND
port 17 nsew ground default
rlabel metal5 s 1056 18316 26360 18636 6 VGND
port 17 nsew ground default
rlabel metal5 s 1056 12060 26360 12380 6 VGND
port 17 nsew ground default
rlabel metal5 s 1056 5804 26360 6124 6 VGND
port 17 nsew ground default
rlabel metal4 s 23661 2128 23981 27248 6 VGND
port 17 nsew ground default
rlabel metal4 s 17359 2128 17679 27248 6 VGND
port 17 nsew ground default
rlabel metal4 s 11057 2128 11377 27248 6 VGND
port 17 nsew ground default
rlabel metal4 s 4755 2128 5075 27248 6 VGND
port 17 nsew ground default
rlabel metal5 s 1056 23912 26360 24232 6 VPWR
port 18 nsew power default
rlabel metal5 s 1056 17656 26360 17976 6 VPWR
port 18 nsew power default
rlabel metal5 s 1056 11400 26360 11720 6 VPWR
port 18 nsew power default
rlabel metal5 s 1056 5144 26360 5464 6 VPWR
port 18 nsew power default
rlabel metal4 s 23001 2128 23321 27248 6 VPWR
port 18 nsew power default
rlabel metal4 s 16699 2128 17019 27248 6 VPWR
port 18 nsew power default
rlabel metal4 s 10397 2128 10717 27248 6 VPWR
port 18 nsew power default
rlabel metal4 s 4095 2128 4415 27248 6 VPWR
port 18 nsew power default
rlabel metal2 s 3882 0 3938 800 6 d1[0]
port 19 nsew
rlabel metal2 s 7746 0 7802 800 6 d1[1]
port 20 nsew
rlabel metal3 s 26681 4088 27481 4208 6 d1[2]
port 21 nsew
rlabel metal2 s 11610 0 11666 800 6 d1[3]
port 22 nsew
rlabel metal3 s 26681 21088 27481 21208 6 d1[4]
port 23 nsew
rlabel metal3 s 26681 25168 27481 25288 6 d1[5]
port 24 nsew
rlabel metal3 s 0 21088 800 21208 6 d2[0]
port 25 nsew
rlabel metal2 s 15474 28825 15530 29625 6 d2[1]
port 26 nsew
rlabel metal2 s 15474 0 15530 800 6 d2[2]
port 27 nsew
rlabel metal3 s 0 16328 800 16448 6 d2[3]
port 28 nsew
rlabel metal3 s 0 29248 800 29368 6 d2[4]
port 29 nsew
rlabel metal3 s 26681 12928 27481 13048 6 d2[5]
port 30 nsew
<< properties >>
string FIXED_BBOX 0 0 27481 29625
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2550064
string GDS_FILE /foss/designs/Synopsys/rtl5/openlane/Top/runs/test/results/signoff/Top.magic.gds
string GDS_START 508732
<< end >>

